`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qunFSkib7n0pgeakP4LCWJE5jcHSbUz30lOfToEsce1YHIl3YHwdqepPzHpnZ3PvJKKRBMF8ojFD
vah/EYUUnw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u4A1x0hqeapczE304Kx6O5EB+pElcWUlZORw8+UCyiozw1c9B9LB90YajImJ2A0DlhalCDZKEpTM
4PqurpsO0E0wVqwivdhNlYk0CtJuzbdpwFgzzMYteezvNKmxFnysSuqtBbo3iCqqkfNg+XQhJV7a
km1poYQEpY8BUDDFiTQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YcJyO/Eu0gyaHauo15HYRH1ssrbLSxq6veJo3jpTcilroOrG/ddFzNT3vNRWpcJBqUoKhN57sMAI
CDZ/st/d5RtMMPeeD9nX2+8GlgHiPfI8CVC/LmR9QhfxTPDSlMPZD+z4wFt6C7hnCa5OWxk5xcZW
HSRd4e1/jFwVhR3Au18TkpGbxsjhAyAnxWKFzu7yik91usG20+8lGTf173Bqy7A9DNQbopVSnrIX
i6xq2z6WJWiRgy/ivGzDEBE4eNm8yYpqoHbwf1eWaV3WNzbZBJ4Iuev4kLAxd5yJBvXL5bibJxbc
YQYHGWmPnyFnUrVo336q69G4/n/yaF7cGnr8SQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sQ3wHEXp+cnbfkiFvXtvD86D/3BWsKuZrbXSmWFRkROkj3LgjhhT6nFQW7OAFuGshsGOYX6HEEg+
k7uAu13uF+V2Td+c9CzxTRcT6Z7DNPZTQYDC2bktvB4yZ3a5HRmYvU/FBicspJfBZXU85tJnnHJ3
RjfmomeTGhtYKsqGn86CiLQn8hSimhB1yJW5sQ6/spxX4HBPSxuX2tQvKsygBx3THQK5sqlhk9Ox
+BqvttrLEImFGI5zFYyA5fa4Q8cJI5VjluKfzg5Cj3o2i0pLoP9XQy5NGZ7+EpUFUhQrBGbO6wz1
abLd7n/6tH3pMe6POU1x21y3bR+xirUSb1UuvA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G8nHzRBECowG08ayR21oizBaAVjYVPcsO/lg4rJsg/GX0ozUypOYVsS/m0GjVcG/h4L5743BhhUr
+h5rKaWDy9DchVyJ+REYTF4n17E4i3GsE1iB62JWriabOt/eZlxUUCjIwRym5ITrNNQAZzLloBvX
mPHdd/f35ZKADAXiRsXbPFN+ty1TPP5eOPlIF1QxV9tSi0BaMkYAVhz+BWbNY9e5Hi3q95WalIw+
7WN7stPRbfivZkGdpyQxVf0JXrWTJQOB3KG2fPkxRelr0Y8JG/tNYIiVyLHWS92ifUcY+15a06m4
NxBs0Rt3+mdvfBnMAOT+i95hsObI7gnVssBkwQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q8YvGBB5FcCjvGWlxDR6zNBRkRjt37zH8JDr1YfHDZ8t0SK6j/CBuEQkwiwMljROjl3qJrZ2LlPI
B/EI2DxTcToZzIuzglr7mdGsOzlbSUeFUR9IfIbC7QQEyFEx+cfECl2P9j8F9HK0oVbmo3cDNLhm
PCTgaF+o8335VDn/d6Q=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y0CjutCiylerP6EXZRZtpTSZnZyg969knomUOesut6JK0hiPq40bKwkzDIg1ug7GIreqF9jr163e
/EAUAiUCRG7/Oth16vE3rYIlY9wVdEIjVmQNNY4TCv1CcX97PIHytAWg4o02cp224zCf1Ft8uuyU
2LgDW7ZGpWm5w2DEw2VK+FCuN+rcaL163uReqBAXJKVPhXBIL+2EaZZQxv4qNb/kJs56wxkEbFTF
LoMRpGs2apkDzvqMmdOWGYfpzbCcqtgka2kX9ZxkJXqx+UCUh4+XBQDWlxKw/2EdbblEZDxQK5XM
ybk3gloL69av2xTblJSct+pDhWgMW5jNUX302A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64160)
`protect data_block
zE8MUssKf5yD9FJXR7BT8T+tcCZjkj3KuCQT0/I166nFVsFYDUhj2d0v3ogREiriT9rVyBbDoI4s
Uby2UKEhm5V28Q5xIGpP/3tvo0eH1K1RfNU64MKTmuwBX4YAG6G1/R96uzNmmqDgXoh0VX2wkvM3
jVtjb+wTrQYgt4qfw8GgSQor48uNCWf2gGLZfPHDy/wsaCY3LQ6hRkJmkLnyj8JSNmjfcrlyVQSu
bOiXljVENylLSguAWlTiVhv7N7iganoVWi5iN1MHZQSCNx2SZx9iZfmpIJBleA27ZRDHygYCvNO8
Axa92w4ggE4DjYtIU/vOAF9gWtXJM5Y7LRpGfHmBOe27ojM1XWFvig/dXOHSwXuYH9G2vtVB6Wnr
GBBngpxeXv+zeBZlhua4HMVIkBqJwIZPxDxWBbw7Qzzu8YYsDeVaRoq2dZym8vf7gd0jg1s6rwdF
/CvfeKxOueg3VEi+xB9FfO70ESRRm2SCb2GW9UTzkyKiUCiNu2PmTvpDUC1RWEdpZs3s6BrObBHC
Z39RYqZs7gGud7AA8jkWxIZMYg7BjYJuZhyr8k9zPS8QyC+wjm+lcE+1fdF51oSKimcN7xJAgFkO
McKyEiBUVY+lW7lEQ7Un5nczEfpx3q20wgfj8cF+q5YFPypDDlUe6yqGFI2sAElOeP8iWs2LBjlA
BkFLwddG/ra18EOCzVnnlXKUWaVrg2r/lzmTESUhLZGpAxD6tnTvXKwvvyqs/xbEw7HcYPSD+/Jt
lSm+QPKlx5T/AXP2/jNTMh6AQVMhRoAP1mqde9mmSjgQcK2sSaowd+I8rzBKgIqN2S3pKU56oeVU
OauPjowGJcEC8Xjdg+U/hJF1eQ0et9R6RoJCbONxpBaDJrnDs0Fse9z6T+liEiC3VrVcTAUSVaqe
GwZ3II88DbmjQXNdYzEVDOQR43NuExyplgiW3LpJR+1uP2bfE2bN5upLALZPvyCxwIAvfA1FAxp9
FXssA7ihXXg3bn1b2UlSMeXeIQkr0sjlPLGHzu2WnMr+nSqiYUXXIrUMtzfWixC9uxpqiEOP0dyh
c550B24lOFrvsqKwLPrk34Lw8KAOPav/htaq0WmhWukzT78lcdoLzHuKKKl63AONi/IF+PS5BgRG
fz8NK38RnNeCiWNJpu3I8DI04mQk3aR2F/fcQHUJS8wJ4jlNNRrUMIzRb0uSNoG1vjfeyZDO4QAW
vZ1o122/Fwf1yzOWbWC6XNhmtRln+YN0oJMcrCtxkKUB42KBkoCzJr638Li+3BvTkn0z2jri7YBi
9WWHjBDmYWmZ9L34u2pWWh8yamwr72bZRJbJGT2C7Jn8IBM6n5MMyEP9ALtuwW1RDXM3EPjq3h4A
/ydTufb/LlLdwvPli7J+3vnhqUqGXmdmabIM2cRl/8nvKrCNV7a6hgMxZ7Nv6K1cNEOWLjsHAZqC
1oUMIgASyYMMQZhskp/Cy+ugkfIhFjC4qzGL/lzTLk13Mu3PDznIZCpPe/sXNO4dfpDsZtpV/B6w
vtZZrS42jd2Mz/TgQHtaW6nOw2jfr0W++/LAY8VamYKH/OUl00J8id2UeLbLNympJ2K+GEDYHJJL
9VUusVZydYHFNVXcgN4ipHEBig4ye12KYEnP7fxHLJhkjMhrBb3vxRAJV7j89aL7lik8IOarLApZ
perr33xHo1cMlf9Tg2trBqwZy7S6D5MJnSSV8WNEE52j4DZ0rS5gprexg/KNE3ORqBvqgHckNIAe
e+Aoqh6zOM5O5E2PDeE4/KFuXVJmropzCKmC9jrXiwBLHYCW7Y2agKd2IUNnxbgRuEd9WzQYDjgp
e0Csb4zDucwIsaEZTEoLBC2ABmd6DwpIq2MBmhQMRYsKmZaLec1XZJkFBW/NaB818pybxq62vZ0c
qoyk/qgMps9rF0BvzSR+o+u8Belv+hxNCSo7xLLm8OT/bO/9Jd4LiBdLNH65xfbTlj0yg1gBvq0M
ht7Uxqfiiwht9i/062p9wznUlRHLKyzqhW8r7ywK6baUZN9PjXhxy6I8iEhgkj/x5wGduihu6Mg9
3JQOXxJcl638xs/FuITjDnQo6kNZF2UD+YkNKjPEGf05U6l2z3X5G4oc3irxw61Zjuh3wdq64lvV
2vH1sOlpjnlJ98WU4fnS1R6vA9tX2k1qAWQbzhVMrGReEcyvui6LGRYXRk9DylRqGSxI8kpsmHH7
zp6X+uXaKSSxYMShfKUE5UhgfudSPFg8VTJmXFq/jDBbSDbuFXBVF07yXXq3o0vzXa7EM9JwHlip
f1nUYc7tIvtH2P2811Ldn1jlvmZXytn7NHA9+WbBwOf62WcsDXvbtYjgZC+zSbEF4jCan9Pnyh6t
DjIOjv7IzA4hP9VW5dPxkchm2nJ1UyHY20SWKUDrC/nF9WfVdk8hzZ2le4zOyOZnMyWjwqjKlK9r
9D80OYC62fxk+LNEcIcsDP02v84osPp7aHEeajgFFy+WrRrP30Lwfeo5ahDWTmB+/aFfvcfO9ypF
YR+8L/6zR57hOpPkn5MUb2YxY80aQdnEqaRAB46rndYtlBpDsQWZvEDshKX3k6VI9Jq9yCHdMc/M
mgjL/G0h7ywtzRXaOQY7+sppJKYo2lQGum1b3XveoDWIG/+8KCc7t7NJRCvF8/GCsr5UDVcGfdWu
cKC2bVj+ZK/N8GYIkV2o6c2N1gC2pHsNYq5VXWmGEk6TDxGmKT0e+bihGH5cOhoZwaeI2y21o2mt
qn1HhvhHiZ7i6M4b1fmL4Cr/Zz6tVmYevWgnUUf+ztk0VH5Qa69R+rAxcKAswBT5dciJDqmh8J7Y
iX1qehAncEZJ4JR4f8V3uZN8bWNB8grWBmu3ZtUd5xkK5VgQmuWRtVhnAO2dl//XYW4/Uorcg5+g
vf+abDJ6ya1MblGeH/YPUp0HoRBpGnf4Y1ALJXsEgINEOKOWmZAN2Mlbg+chrJT2W7Og+WiHGOaP
Vp1LSecTbg35OPzKEET74GIKcLjXDq72FMdpHyPfe68O34m+GTlelxdpJmUyzx+YZhLYU37yCpXb
hNsm15D9CAMS1NQhIE3m1N9oEcrVio5RzIWDpS9QVhPoaSLPhHve21CSbrWvSsH5jNSCMGMtJ/mM
BwCiP7FZhoydoNKcsrRRKMKPV2h0V0CmGookgsv2p0VZrK6oZvR5jTMWhqo5IomFMeblf/2Wj3Qq
ojUFNxPsrIuZ4yAhwvMtp6ErId2w6gKCxilzcKneGDa+j3TZJQG/3mdal/iRYUIjrgxsPk3segQ0
9y9jNyoULWWBjb6cDT5cDMlRAcFyg4FF6n3kTLXqbpvDkClUwODokEXci/uk1y4+h0QzhvPtfPMe
q3NR9I9r7AoC/3xu00m6eTZuX8cofz3ZQ/wsqCqF6b+UR/Tkso6/CyhxIXFECk3V6uHMomy/kktY
gkHP8bWVHR/VmJnXR2F1iFzKJ1CnrTc4AeK294hpyiyL+gzqPiLg4UzwhL5udggSPxEQX0Banxf0
F7TlmJ6is7fSQEbk5j/zicHwqd6sCuYr1upJCYqzzlsMKNpP1RJbE5wwuM1uHJlp9uDuyEBYUzjM
wyW33u0nTupPlnvd3mWBVLLFyKhUtBh/2BEgRc9/ZBOQms3TV61Xl70RUG4Me0dpFFDghueW+u0+
us7rBLoiuty5Gz6a2x03CbdCu046n2UvkiFOtmL72dQdQ0JmoBX6omkkG8TfHd26hAV0SZRmte+w
F81ch/Gy0xA2wk69ZcxZmewUDpnvhl9QWVvXnzgd2M44Kx6XREeZ1kGs05MVJAJbjg5qMW5LMy6A
Jkt+940CI3q8tjh8IbFbNr/rZ2WA2DYXSHAfNJ6mjmvUTLcaOHEjgRwUE04QpuGrGJ3lw5scb6s9
SWQ7ERagJTlualdW++P8YkRNaO4SHJkrmxkP7FdLe9XgNwsXzOKB6vMre8yTP31ozFwiy/+m7M+U
sU3mNkMorMAiQpGT+LIsL2J2c1VSplr/N0OW5xJdnX2H3LIbllV4GAvQaSSqHDsGzX/ktNMNf10t
aoSNhJFxKqAEV2Leu86A1FeMf5/Tzl9Da3Oi581fSZv6wIuvGYTWiLnU/mdB6Zoewv9gcPTtnkbx
dxjEDdFX+o9NzRaj7/cG/WuT3rt2WJ9HXxO31ZQ2nav3LV/CaxRyd5e7pBPCsu3OfGXX7pRxvSYr
uahDargxlel/8dG+x0rrAJ+wmFX5odDQojRH64q2vARWrNG04rKjnGTOwrPOu8XHrT+J2PNrim4A
td7FY4TTg5EPCVZWWbOSCRw8BFlCKSHP+pN22JaJEHUglKaARiqlMhWPga3RK27L6/CGPOsy37fs
GXDHS5BmNTZ6OduUCgvhQGNB921sGAcSz7eiTpDpKZgP6n1GzSKSb1X7AtNWw+HhCaUDgdcmWxIU
wWSsNLouhqdDnuBBO8JmyQt0qH9QG+KhDy/s5ALrInhb9epF6gO9rlnjiWjiRwt9AqFD5HbRd79b
SK0xYgZCsycOrI4Zs3QGZPzVqSDOALBCttVEzk191ukeqb7r2NfkBICRjvD4n7Ga8V9Y4+QDlMR7
7qAN6M1xurEpvKOiHeA0tUmFDdAVnzS0Nuhd9Qo9C8UrZEJvxfSMagxSUnZMeVm+YfkAAo2xVXd8
GneZGDQHAr0h0YQEuDw8rvaIkQOjEqFTZkT+7DhnEOQ+PMacl4RRX35Uzp+srYrj0UsHnadGExEk
zmFD/IzwtKZ6XQjDbiaPqaqW5mRbiiG2zFap4a6BHJ/5pW3X7cjHU9L76BKLNukRxiNdmwCKBqfH
5d92Lfdv0QJQcY0k9q/Bt6EFJpexCCCAZ7ZqV5Gk091dZscQ3rUs+6oKRUDKWQsjRJNBY32qndXC
YjMOtZMmPuv75cIlEpVGOBJSiycp/QnwJ1etTuuaBXRvQdfIkgoVkDsZGU5qsGpxrj2g23nNZs6O
4dWnUvgpsqctxVqzF2udokO3lshKWtrr53URy+AsGQWXo6bQ3Kzzh0eKE+0hyy394P2mtEqPfXhR
5FgGBzhsQyTJPX5Y6gRTDmlpRwI8J6nlx8TS3PRvy1KqRWoy+5Op06pdByRv5FDifLvQWkulrUVd
bgmO3pKeCXQ1b0cJydSWFlVtq3FyEw3INZH6Btzi0/oaPzNX/ZgAZZOcpdrXviRupHiAyd2hK7eP
hmYfGFdQr9bWFKRTyXk68u6+5hCk/pTa9DOc+v/EQRrsTX6XnniBPuc3HRgkTxuEiCqLo1OjQoZZ
xUdxoIEPGfesOgTpQoK0kNRBE+89x0rRpmYbML9QtSWJw3sPZW+LyyKqKdvhcsvhey7hjAfkrvil
Zz1YZ7Ry63xqKHykCTJEz/2mGA+lPdhWWWldCvEabjlddfNoyPr32HlgFXAdbHXxrNssxR/lNEQ6
Preg+XO/J9dwQX3F7r9YkzPlrKpbZ2w+BFiUsS7g7nGvys76e7qEAxYvwMbptjGd10Y02XSKB1Bv
co4ePHjIX5hFGVzeDXNHfNTAMqYECjIQHVxYk6mf/HbKcBHU+x69BL7mZ0InPWSrW30cb35T17Av
E5evsFCOlhuwHnuyoYmiFgszV1BzucQeiPP9wZAmgzc4lQPb6hApuJav1SnMXTqXof/WcGGu/+80
yac1HjeEJUuJcn0Qkcx+RQ86OlhZQCR/OUHn8YIZV3SesjIe/5S+a/RArq0TYycWAz2oxQ2uA4mL
vNm+A1ZMCnVLqWtcAw1LvjSrFtojdy+S/HyMcxsu7MCY3dihdIyBWV88fllO2AxhrAFiXSNN8WCO
7tyznoH6MGwIc5X0Ev0nzO6EiEpvoN++8o5GOjR1rWqGjyatLa5+Za6+kKsCBy1mJ5vSIuEzNKQY
/Os1zbJU/vEiIj4r1qW+1HcrH4Y6W905pORc+szOhU9Mv+NinG0D5FcswbGyEjnkpDbYM6WE//+t
HW1Db8PYxfeTah6x50AxT5vGxXS/YEiJMsrpF0aGAmKlUuVGHqsRLK/emSyVXVLpNzj7a4fy+dC/
ra5NBDLW9EpaHrsTHf+YHUMw3KRgIShqIRa6aUyZbwqFeiIeCUGY9bYHJSsof0Z5vuUcQ6RSSc0N
gYtA7S1iAV/SFlZGVVTrS7qXiAMm0jKSnfQHWJ1DmdE2Z4v64L5SjyOfDu36+BglMnzhefyJ9nnJ
75MDUSa4VkAVc3NPXwg8e5hZbO0Re50J0KbFkyon5yviZldmiaKV3YkK2pjf6llIby6MoHFTyJD4
g3lybpJUjKBjPdE1nsRf3UGAHMWDBwVbTAE8yvaGbtID2lrbS2E2zYLwRXxqVuZXma1AhmQtap3L
rfqd9q4tYr2HSPnGF2zkBO2c/SFgKBRnThjnVZq2Vpnuo230rQn610LTBRfbRtDAoo+/Dzr7NHwj
S47W8iIYq5fXHvP8WuXe2OwYMHaHsGk2MI1lxIVZXOYV6LjsRBZThdeQ7TipRCv3/TmgxnQX8Jwa
tUvST9GHQdBFgjse+ZlLwhzs5mll8C0G9Qv4GC1hFLS5nw2tXl+zKMq7lJoPYqzIJM+s0IpkIzX3
tykeuCC8gYYHyx9gPiVZjiAkw9Ukk9MChzT95E5cW+VOrb2tdWjcWN44jj9ecZHI6tVHh/x0JTvW
ghRmlU60AFvAKsgPDA7ZiR3Dz4elVCyJqwkmVEGKVL7wcw2KZdMmLxlVVwEwbxWFEfrenEjNGDmI
XQ3CxkbzEQ1fFanzw+asYX+i1SuAxKSFp5cYTkchPOfPd/8WVc+SZqWiJ3y/2gjitVt79EQcQYbr
b83H6NYVUrLq8sJRPCZn4m0vM5Hixk0T6a2X871aZgzTZO+FprrqDrFvnNacacA6yHvQFHKzlIA9
fV7Phskxsc+6RAAPuqz8RUtplzNRMqDPLMFO5+5YWzgtjgGyBfOalxjHYiStXaI8Vlvbw9hdH2Yd
rDQvZj6oOZrif30tXU5LMYJHyaRa9FYKZR+2GDql7cd+wRtZ3619PTfY3Uu/gVLJBjxpmcRSfR1T
5RRHNnG1ditdDyRjgSzFedBvBm6nCuoIikthnbxM34nmdn4SaacEg7w9WizNDKE34QqUN2PCkrMY
1S2EgIzh0tD8FWbVM1l6I28j9PJ0OqkpaPz4xvgLsXOBnrBDIa+S/tLxVD688IY4YhHImRE4bMTj
OUwgNi5B81lYz7Wx5tGq0iif242cDi/oPNQxuZx/jGiXkYD3rZp8aIgQypn6viCGL5bKlh9nkg03
PDz1EdlUYi9gS+TMe3/c0k6rFeQzQwMp5xHQUuSM5bfKyBHrJ3ehO51xJbxfkG6qeVgLsMHqOmHm
hTb9K2O3YOkZ+fKdjzM7S+Ktu40DHMatFzewrxMTGjRb76rxFPPg4xL/+5S+Sv3kZy2dQcfKsxS6
+F+lAkQTYB9vjMorLTejPX2juOQUAm+B6iBvjUVhNBUARB+HbqVHieihfbNYyT+ZG0p8rYiswlW7
lGNc2xM9MOe2jby6jV+DvGR2Szguvf5NL5fTXgk+k8N/GD6UgGznd+W7TvdJUtSdGZhZA/MVWOvn
+kUvISLE5QufM7uYro6z2r0bx8jfjKB1iNK/J7GhS1iXNM2xBix+otI0QYBh3TAKwseM0nV3NmJu
7JMChHxfxz6/zlNs5YabhkR2Nj5lO0wEQTwQ6E6R7jPv2OvB0+3qAspxaJFxc6nRZWYcBeH2IyEk
bIBiY3XVgBgG0Uvno2MDd7o6mxI2Z0H/NJgPIip4wbvoY3ekQe61jmuPAzTczIo5u4FOE8eWCbNr
DiLxN4nT7FuuudvRRBynCpKm4sF8wC4iKFTzKwCZqnkVks8nkX/4XIbmrkzt/WOpsGPXB7Sj1KTZ
6suzaNbwYlUhRTjSGaWrVbAWrgkV/hUG+pDNp/6jFkFzWNZYzNxaAIFVTf/DX3sOrzov+SKJxkBB
0sXOIDWu90mBReue54QMjLjsDphs96QEk7yPoHmAX0yv4qyJw1tl7v80SxXWvM4Gf9mYkKzyoaqD
ybbj2JWPx3UAAx2RfAX1e+rOlfUnR5Il2bWZrj6RO6uMK6q/jfrbxfDE+T6V5HUZyI8BYDYcy5ep
tfOS4XkEQedQ/c6cv6/yeNBqRTb6Xppnvudp5Hmdh0qJJGHokMQF2RkHhBwCg9R1suorJGkbvGjw
yZyEuzYxXYgE/rjQR5qks1pMrwZTU+n2Y1eJBChZ5OVz68MDMibpCaYdPR19pmwR0zfQG3MmTL+y
+l70rpKgkErVv+wILs/WfGSvV+4ZiW/AoYBYSBgo6svKpj8M94ZdS/F+p6/I/Z/sOouzEEonP3OC
Bas8g+FL6fXOg1ea99I1B3j54YMu9kVl65yJ1hPaDo/w1or+6pWJXGTchX6TQKufwSBlSPmwsYPI
yY0YIpUG+UT5l4apc5LEJ720fMOiwSmw2pzTgfFzDMpL6goY9xj6gGhR8gTMpMhFuZp9T0n0pugS
wXST3zv1kzL+eCF4nxqjkhYrTQi1FroS09yetOqxvJ7W70sDbo1Gw7YGp+GX+UpDguBLw9HB+2K2
PrGCbxGJRIE/DybQkCk7wp7R+eOA3LvNQsL3FIv/Xbfh93vBLZzYTb+dnd4sUEOzdbcj/1WVlyav
lXYekkKsu3Z1QZ6/J6m3CyF9SaPpUuo2LyBvfgaygkhbG4+QbBbxNjwG5Yo6ZUtCnLcp6Iu0N7lR
Pp1cfoYbBzEimZexN+FGPKUiGuYh5tqonOA/whMN5HnHAjYecZgenlhkACJR1KoXOGGJ5VTSNV7H
3nhZnAkK2CZIycfbOmj/60olkt4xLAZ35lMlgNADAvV4kihTb4XSF+WhDL59zJchlPWegGhtdxOJ
rx6EKQxSfu9ifLB2BJV7tDz2uXutnvc4rDdfXBbGYzlkPMOSEBtaAU2cTxGNrktCC4dnee1U7Hi9
hIb3w5rl3Pdm01Yjn2wO2h0rIznwyrOH03rcvNlxgx32UETLF3oTOgJk+Of1hV4q2+YUTfFe1koL
vn/xe3I/+joQTynPy2IrHCZvfWxkmHamCOMb38BZPSULxl+Qv+5ZHq5vN7CqM/Y7xDZ553J4MywV
ReUv4O2jGK9seV3BVAXL31IEujmFLq2gWOFV6LAzoawFfbDY1hWLit5kllCtNxk7QDg8IpD6/fr2
iSohTv0efPqVePDLvmIRL6dSNwmIW2jpMTn1s607tc8pUoO+mV/RaesPCdLnYY/WJWP9I8U76XVw
GV5UPBd01L914Gs4NM6y6ZRhZWoHGihtIVGNNLosltkQAAO5Zc4HuRk4L2IM0JDSKF9nnGqhzdZC
VrFywwRZPVpZwo8z0kMVu86GGzN279UFudX3xvyLQYueQvIuZG31TnQMh5W7wvm2kjd0EbkBIiKV
uc9iTkn3bmlHIhxZURuvQiAgsHQuBQujlSGMLqHVGQWnwFnu+xWHXlCvFiO087KJxnxcYjPd+u+P
YxJkERHozU3qijw3oXFSad0jQwaUAu9v1Jx6mfASXUieGNI3RUC4lxwQrecaAfW8B9vLtVqbTf2x
ziFwAQpWvv9QaqAch1AySee+GuwELiIcHbwpQaCMrdRuOgTgKx0jGrRHyVc5CY2ixMxzpjaKR+r0
v1evR84Z8y6b41UGlAS0HcPG29TJADrr0NztK2qm6Zkgqw+As01KQSQkwymz7A58VcvLFPeQ3+r/
Mx8SiW0I5jz1vK4ed/NByUIvCySJPOGBSpTAbinjh4GgKRxajvC56hFE1lD7OzG+aksWlTTOxyik
Uaxkdmf5sq79NahlwQIka0y/vVKrVELymAS3WXNkq/MKircFGpiKiQrhTQVre2vbfHMzAiZPSQcy
5uarMfThrQwv8hph/42EhBaDs7uvJU+/REYvpL7+scKckV6c3GiOVnK+8sWEnI5qSI20CgjbEj+7
9nwevUSZDOCNtXAduMtGOzICbaGXdAAh6ysaziMq9rKe5VlXkAkx3Drxh2PXcbz/m6RakZT1lZNr
YRRSM8YpI+KCeSzffH/+PJZfJH+IYVs82gs0ynJ03+OyJnnkcPVCeXb7OaFm4+oGt56BGSxVZTc8
7kqaYEDF8tgqE2qbD8nmhVdBeCuHAnPzxNkp3ZpE06CmnPPSZcTHIx9okNvyM1YVHcyGozyhKpMZ
HgUZcmTUr0HWjzo+o/lH5CPAPq527hI0Xk00WeP84ih/KPy2pI3WRKMyAAz4QkJWYS4sGyvN6rDZ
hVKOwJGpfaoQp1ty7Oofh6/R/5a+Hpwzsjq2tHiCDRn/sKCZIcfvJKG49rmSPTaAfB/IcTIQsQa2
ZQioTUf5VAj4CnW0oMMQHc3baI7XP5VTl/lsfw5/YitJIjuA4AsUGO6iWb3bTUQom7Q2vTPTv3Ff
celR2rQItZqvDhhFIPkAvBDs4PPu5Iymnc919YaELll+BU4B4Scw0YSlrOIYTw2r29keSxG4gnLZ
GSn8tQj5SvJg/xmaWrGpgVZR+lOFc+Mvj2anpX7S2uwUYaRzxO+j4qWJtPgxQ363HMz/y6ZVs8kN
nqPNMe940zuq/Dv9fxjppFg3wq2hV5ot6nqTZfNpM4qJo+3cBZBETlbNj76p9zCPRoqFWmf0xQPQ
UY71gMcIt9+bg7i5n23e7F58UZ+TVUoiLkRaRa2o3Oa6oIQwKTN4vyaH/v8wld8i41g8NfCKa+g8
R4C91zXgNMC0+1oeJcijke8NGfMzBbLEbe8KY7uvjSSJjHg58NGDqX8IMMFQbd8kZMqe3BTnzary
+Y6wZP6335xxGLyTGlKFwcWV/W0veDke0J3Cqp5R8ezKbfJlPH4grFzCFz68o62eOOR7eDhxTCRW
FKCPpzR3X+mHOsXddaPJxWTa7oktPI7U674HGZ1EBJBoaJTgK7FglU/qjjvPA3kQ2qi4e3WoQ/gb
SCoKZVOzMBOLrAEHiL8CAd4DPKL3WrX+8Dw8QHMzt1gWUC3nnsIlNN1r33cRhYhaFqkVJIO+xBQU
u4WZwIP7Tr7EJpqcFj3+w5jErCz/noGsDH8Qz2woxULQ3FRe/Udl9MNaC6qkiP/QJMgoUVaIBguA
Lk0oS6DMFIHJTmjYEK/h5A6cnHmrEu01E9kVqnpGZAAv6IH6ORkkAHwaRP2Ur7BkSiw50XKLswky
8f/B3hMmwxsnBRc7CRiRfA8UJCim/5j2+W+RnzEmY7jIu2ZslOtZh+k5JAQ046beQS0kEYY4Fsxo
QF0pjLdlTQuIfWNdRuR3RiK7L+gTyEVP09FCUqUp0BmlMGXa+1gEelbuKspJmC2EMCCDxE05760m
5SyRekBSNNkgZTOKUJFiFM5B2AeSY2V0rJYIpP2/eZHFLmRUjSqzksThr4oVnMxlGdgjZiXah9KT
xaP8G/dnCfxZFEKWBanpG3I69WdLovcX9P/n2gTOA2fjcY0U4H67J4RmhPooej7OBW1PfEOMQoOk
wY8qmI83x56HN53WvM+d8yD45q1lqLDz9HhiHys9CdOK0Tzm6p5zMv4nknu4co1k2prgeLgrnpv/
8xlnzv5J/wfEKalL0xnYR6yDGJHQMD66ck/BpfPubinjtaSLmBJNNGAEZtUOUmFwf0y51WeCFda4
Ovp6HLVea5h1dVHDN28IkyXAnBsb4Fy1ClyWIzcV9POoUDxz193aiBAa8HUbsLg9lm1FF81qmdEk
V2l36cKEcJkD5TzMIMk+kfXeZdWElVL7qV82UH1t/s4L0xSNKYsPjtE8yzBrn+Se2LvXm1I302bh
4ainpe1STflH7qz9+QG4dMQ6WeqWE1jMAtVyW8ctm1Mti+6kLj6xiWes6xFZ/bDvnKyctFJuuUCg
piu+sur9LY+ZOHD849hWSM4uK0JPMq+vsMDPchEUPki4KFBTEd0ibqFjvWECxXH1Aseq0RdxKGFB
5nkrK2AaFXcPUIlxAYZDpa7vx9j+fW15FibR4Dkx6naUCXfo/FYKngwCQ1ZNaOryGMHulG+xqpOg
V1Em+rYrvfWTdepiCjAHrFvDfueiJJPAxfOdh2i0vR0vSWN6ZuXW0rkJPPIuvSLkWY9KHxJI17mT
FrwWhY5AqxU665b1WWtmVEPJ/2TWqZMAwGorrgYYUdjoJuS5oNGWwG7UPZs8VwAJGEzBIagr6u0Q
iLv3xv5jbJU8S/B1z/WCWNh5ywlksVSBLhqNRMVLP652mWqm2tw3bzVzGkrHn0/q+dfKGyX4eSWT
55bJ3ghoqD8PUExWxRxbSHRYsyhcqqbgH49O2gxwyKLGfAGHepHh2L1IS+9wju/hXe71TYLQwZnl
BZfqfB6kDIXW8rtR42MHYQlh8E3S+Pg6jw5t8nGKP9jXO75Rnj7nl4NSmO10+D6q1B2vTA0dLhx8
04pZt/vV/L4hSpM3lqTNlOvS8vXLHpfqesng4alsZttmgQ06Ag6xCmH5ZI5tVtgcy6zRxa1Zl9u5
JZb34/rs3Def56IUaQpqO0HLdKp71n8TqEpNQtoeZhQLY25vOdlpeAnR6URhRhD5dUSgIW3CZnBs
v+gImRalRGPvzCLHWOFNEKy0Aak0PulJD6W3kPaNvE34wuLSC6r+2VRHef6ryy1p6hifSuCLieha
33aLMjRPkvfQ2Q+x66U0zxVviZ8kBIbLSy2cxNEJp8eKYQldAacogEvMq93+QMBwtriBTd2Yy1zD
I+2rgUAL3yS5OA+Z7tqm07vqAwN/IXLYfXeDmMUZYXFT9LDBZAZdj+GMqxPFIECaw/ZkYNj5f9US
MbWUqY77YmHSBDU/GR65xFYh5xyqGl1L73rxntgEepD97HPAsJxmOsHytbuy9ZDcLhxg+FEe0lx1
S9tgaLJ0JWRxTIc7MRx16YVBYKA+AH9/xlTPgKuK/Tps8eUuAnRdxQdOSWqZmIOcpyQ5m5omkHF7
bR2XgZ5FRcGsHo2pd+LJQSVyOKKGkSwoZrMuMIFmhAF1XlifK1iWHGTVIJoccmYK9V9zP9a0EpL1
dj3t9bXn4qS1Mk+e37QCSVxeKAzHRwJJyAUFgTElj94VC0NfpLrR3X8czEdDs8p0rj1/iK8t+F8n
Gkqh9J42JkD4uPYC8p0bIkt0TEi1qWRj9DKe3FsgQKunAEIWw9EuGxnyFHPV372Qj+0DSqM4EazL
Su0qmHCjkx07/BlCmIYwygNfV/8VrJBBnwWEIvcZNpZKFehBqVk8VKBNkp9Fp9xe39ye6Zm0lSVd
50mWWtSN9ZrjwLZQNMXcuYt0TCKGo6defxla2H3khXFagP6ktxHTJB3x55wUHN2BwlBZPyURDqEE
FdP5TXy3p2JO72hzAa1w8Y0x/E2Dwm35+1xA52Ya9uhp54Hz+ERbk7qnR+ZYtk8o//z3GjhexKGL
vDdMyydF/Zwxm945UncYqhJrx9YOgqvqsgaUYgiXUDrn/XbUnAWwBYCRDxc+r54qHX4gAx144Sy8
EIYKrTyVeRt8n6w25XP89UcnEon/mVew373KT37irgJCJa/KBT8LucP55XNxeqcFTO9dqZlmOXUD
Ppi93q/a4ujnuo8CIEvZBhIsYZZMcv4fMTjmQRtyJ6Yaj20vLtX4oy5nFR8LggGxqY+Jo6lt2edU
nmexgOJ08Y2BWWKtD1sZXrIdcvYlY+w3CKepDty/Hvl2q0vv+L5DRohtW58odKURT1HPnNNuZTAs
zf365DPgEeNHw7J9cHonwEuHA6WSy6L5drekDDMA2F/avaIR7sGoyN7ySdiGAcVJ72bHB8AMcYgc
tNZmkC0dLDscutsTeCC4CwyQFM9qQL27owvJ8LuJMXAuS81SAFYfqc1nUsqs4QeVxrXMTvZuT6qa
ZbmokoOGqbx5w5M/vY2eGFXfGBHPb/1PTkSLS2tpr+eWlFAlX4nH6EkPOcBOL1ZSlo1VRIUT7uAs
XMcooBIMupqp//KEnf/w4m5fvs/iLL9aN4BmAgotJxh3vF1v578QoqloigBEiF7x5wihmjWlmiRi
D2iWFbFb0TegFym0QRDLJjO/yQJpMn7RjVCBajuj0xJkhAiomnACioqQyRnit4fym2QmVjhCSVY7
F0tHrMYOLuKIU0u2Cp/WrBVf+JaXbHc1Z/E3P2Hf4co8L0vi03QyYYMHSBxhchrqLKQLxSHUK+B7
rRNj18VQ94MLSJT5C4BrLIP7ZfjqVvPnGxV0TI28Z8OiKmaeOMteAmemf9Mzxyl7psRLMRFIeHwu
04wxfDTINBR3dFYupZ9nUYwJRwKPohL2m+FH8Tpq9mOXzskd5aM7Z9m/uFqCUwP3euUc9+0yydse
1B6lzBbFXrAVS8hNFthP5J5S9aTpqCJZ+3KFNXhsY+bCXhKDJ75tqf1j0Cm3prFeAutHeWaDw1P3
FWZ6lb59s/wsSiQkA58ZET5TNmd3uZWPhALvj5L+SzxXRM5pSi06vopn5U5pxwkJBbGuS4QLTNol
Itm6hiVoaZhJ+7q4+pGgSfRHtl+F1/A2iM0wF8QhwaVve5We50UrCOr1CZUjopo4BaguGRPKughe
bLgjKlEHYwm2epvorAFfOFyb185NdLCEdbMEmzHaOoomXN7kmVLlO3BMyUXFANF2x50ikhQf8EFo
b6JIycNI4+9GC+75rU3nKkNtND7zlK6mUYeJYq/jEl7VWbnaCjCFGpvClzpcsiu3p7JgAoXuPFag
j4JHA325JEEScQ+BpWif6zJiON3ucpQQOtDr8V7KrpqJxkfjGKqDHsS0oTLQkzV4uuo0hwzqQ5cB
h6fQpvJHXFfdhFzyIuzBWAg315wV8n6WNAWpKeNe/d+MLBY4BRy06hkohBABfbYkAgAnYV1hh+Xo
Mb5pc3T5em5IcGlUp/kfTlKWZTDeQFbIbgOGwAVRwANEGkzqblkAdqQGPBC1m8nVA5cmEHn2Kanf
uLfWs5fniNHfXzVzxwfPdGXcuk3wlAOR/25uiytb/9+3PBy0NX828TxmAOv3jrx6M+/OjYX8ebHO
NZ9yv1UWc8o263NFpsd5Czv6xYt2mx+0QndNIW3sg9xWjboYwgoHRoi5MCpsu0r7n2pDibPMGZRx
IjSGw5xMoN8Xs6g5HUNcJZEmEznx5SptURw3JzuB5nfHV1/F+z3rQD3mj+NjYQJ0hwcm7ES4euBI
FZVEpapaPJFBYdXN73gcjBiTISYNXXUoUGhIeNnKA4LYgNN++m7vB9AEhB+96JnImGkv1c0rgMem
vpfyLgcNfaIgidrfCVmtjo3A7/7SH/QC927yhVvF6Rr1f+BRx5LmrpF1yvny0wOIk57P25a7vxVX
BLDnUtn144KaXVSYT3raKTeGtKrfnaRmQqIivsKu6e3qoDJw0KZJyRf45OFGlHlfDUYBOayB4SFb
VYT+mcEM3ZkeLEi5Yzv2LLJH06Xt67NyQMtWCYM5zIygADzM46HtkeocCs5aUJaC2KgzkmT4735k
3U0PRrMA5TmwTZNm3l6emqIc5pfuEEZdLdOORTmU+hpSq+84pB5xrQuNK+tnEu9gmManWMid63wA
iiw+dLYGYfMCF94Z+vLS6ukIc/3IMI+ZI9Ry8TiGR8DvJlUg/JqLD2eCChqvCBWE8kQ2UIpN+TBD
CdydDz/kPJ3Z3LelHXYnjGd3H3g73oUJZVg/rzqGDPcwVCTe7YTGa4rxXXfpy/B0I+6DOuCb2P2u
jvtOwMfs6fYGWwWUkbhAXz4gvUEWg5qSvdT5+Y6GWhBdDvkrBMqzgGeHLrz0UABH3g67OXGlmfZI
VHWHNCgQ9bDxLNNnnh+g5cf3nVIsCOvIZJ12BOlEESWBhOrxdq4MqjXZIllhnSCXxXYkmJitxYrb
5Pt18JT0eS57vhENjKRdmW+juZ3kWATt54eOBG+U/dpheYeqpG/tmfl8kDogQXqDRX8YVv3Ct8a7
rVrIokIaBImWnbIAwy309jx7dUQNUS8PKUN4WT0AZJzfh6v/QR9NYXhC3XD54vPahSprZNQHiDdS
CeAuTxhkTC37wwts4cPg9eW4lpbjXldRPephinr2G4JzgKuytiiCM9BDBzXHg2B2GUna2arggvc+
rL9OkexQZac/WxIQOPysAb9C+w653dx/ILg4BY7sEqsQNg2qaxaie2ulQwi7fcI5EE4xxlcGY3Oy
8jpWlHyFOzoYbU/Axr+WyoD5oaX4ilTcUGCLdrUMy4Pg+pbaxfQS60IRAEeRzAyc+mzz0fpPX/ZT
uv+tJMdRnGBlQjt800t3xMZA2f89UJrWZkS7gvtomtunbfNuvlF5aGDGXPZ0hGRcVabY9fGGmcE5
rQpThyKslTGgtD7cEc1l0F9xo9ywJ9mH7PHsuTXUqHybEvDh59iu4p0y3RnYJ60KjsCzAofStR+i
HgbliDfhclOHBfhPmoGEq3q9zyRBeddtbIHptg3zyOde7doAkGU5Yc8Ivddbf9ECiii6rnMuVECb
goPjDwX060dT7JaYj+D4uvE9JurD4YPbnvmi9UjKFggBRQ4qAbZDYNxopCUr/LsA6sqaO9Q1ymVx
HcQv6D7jbzwRaQOarO94eU8fPhUIs+jkicmkl0GjckDH9L5DsjEsV3VItYU7QZKy0F3+s4WkBQxx
Zcz6Cp3T60nwQkMO0hm9JLhnVKH3JtVLzWHgYOyAsqFCV3AEDHYb+gsHDcV9FcKXVwcHd0cYMrwO
yvzVpvypVsJvjTNnxOeIihtAhMR449VJMv71/kGBMPkh9JeMfobcTNmUmu6kLzlCfXn+hJDUbuzD
bN+HkoPTBlTNeqTWbGZ8175DmLd6JPhhfjLEWTcF2uBbKvA4baDeX90rZpYoa/6O8x+Id+B7dbNP
uxeNKjh2wVdm6+bziYkfuHHYa6VM4MATrv+Iuiw1mqXNoVcOrd/d4HsM9yFb+KhaChinrOXbBZJg
K9sLpni5afIfNFkm1xx2qOBpMV/c+qlOjGkal6nGIz8x+j7PIM+djtJe93D4uqbS2z/UArQ8S+3U
F0D+BmhyAey3DBnBK5XkjL1mNn4ZXQYP2dFNq1KES24d+ZlouGJX2fCo5NMaPXaQyJsTwGO8e9+N
vswgxfoDTSlH2LkklmAUI+U0xnmc7DfGr54+juk2hJZwllByKXkEDKs1ke/GClXjAo8sgJpwoqfk
tmHBozliUXOVdpjjSzhiQJbgtZzx6H2M12VW5qGTHXwCKD0hRACFvkuJBvlAB5KceuHmLD+X+61y
AneCkNo4CR/zuQV7cOnNLKMozz3i3utQXs7qZHyG0ys24bhaIDRNw3VvVA++zXu8Z8IJ76uPawm4
KiJj44YbRkELZSoqYSeDjf1wdUv15sfjZe3lnb72+hWm3zSooNZhdpJSv+IjwaQBD529Smn7MG7y
TrMjGi0gSgfKgt3a8hJPyQQbVBM/YhiwAncSq523fbpw+Aq+3jbjDwhp6pQ9UAfx49IoMYGKXUQY
UeRUTh10pii48oY4z+h5ZkVZE1n8XalMlvzjfi38fi5PfZKZ+CT/kFuf3QmU13qVIL4FnoMZXW8L
9FixlrN/RkkJtGBDZRiYfID8cfCCrvcP7dlQ9Ivrgixju26TV9oAJfnSgZ2TjA1NspH4rtWGUHd9
ZAkK+075eTOnGxSgfrGwZUDcblv9mHYzV6dk1g00F4RxqSCPww7hf5taWKsgV1ad9VgKOH19po7Q
hcuTTJVKcIFI8MmoX2hbOiXP9xYLjflPZN9cNxtTNOUeqmUX3oEiW66IfbKa+HbWlDwic5eue0Bc
zzqwipyI6QRbZQ1DigBU5r5eCdy7Hx6JHhoAPcpTWqsqwQrqgZftvdXwrM9YtlTrr4+XoRO4bDIC
j5/z613Rpqwrz9E37HE3F9wFW2Mw1xEUMjXhFpr1cFKa73mTZ/tlWmhoN0fgrL94VDe2BZVbisSu
RoZ/Jw34ieAAczUqzJMnBvtBy8tzZn51RXb+wYqdfiamILOQcKhhzcHLg3/CVZylY+7PAxtITQSY
MSTBMyB/82nxwWdPk7MAkHroehvlufs5HP6RX7yZfxxVd0iNYj5Di39z/9qAwuT6vhyits8UUycB
jO+p8P7kLoqNPIWaxgxckiWoQLAU2Jtw1XBXXLTwsxIJYsPqyrZkf7Ou0/qCoI5XNWLbDnTzSXDE
moQYdL+A4PV0ANLWj0aHU9gqlNIOmX7gcvchbgZSkQVr6j5N3cCgc1prXQlLddJriSOri8zZfH38
H8dEtM3TqJGdHCAW8Zm7vwcx1QJDOksPSVkFrsCgmgtL3RViFj3cHbHQ7AI1HLSOjmaKYq3stKwO
6LMSnh66AThWAwdVmm5G1YHrlgo6prR9+erA1vW9kjin7XPG8JfjnvAdHUuPtR+DRRrmB6+LU4z5
oSq2xDeUyIlrRzWbautOqkto+1mxKwDHkYE1oNiCATxeHi8zM6DFcunzxJMvtLNKZ6Z8yEDYenbw
M1+Qfoj25nkKzVWCuq7k7AakAxfL1aXSM77ZM+wodFBUlXFj8vov7TX1+LeslQQrWkYOwTX3tRGl
0r9asukk0TySUjR/VhRQmcO468KFROa/adgHEtk+8EBpcvZMCSxC/gIxYT5v6U/0BQTHcEwXhOJt
TyLiS0kK7ni2NtPliUnxN+Afbm7Cq2yWxbw8hx/TdQTyA1JavrQ37qwuIGOIhKh0MYRR+EDe9E04
6XRLpoAknaaa8yEm1igGhMgCWiT2hzhRTEsUMIhtflN+/PnVoGEyoqck0Ojpoz9nqg6175WxgBUX
kgHcrx5+pWMC9gvBOeVRD4ytiTzROiBnfoUkYnvS/4nk4TbgaMmLJJTzAt9noaLOne2XNAG3ruKj
FMIZtUvYtTpbGe5BmDkxcFuKmSmSZpbvAVKqvfvlRjZ4my52LpYLk08He8QvNRxuCehtYyGjmO8R
n3BhEI9Ni2Z7KRsLuHeai1xwFCPfx7LR91rnhB0lQ7C/p7DydshmK5MxJnN6hK1trRGqibWWj+9j
U2FEhWvoFSs0ZWwChdYR1RgL9Dqk/6iBwXCtaM7F6PDo6Dww5My4YyPt9Tk5H4Y3PwwmCsSE5MbM
yorcxTA1yGb+xZV072M6AEB4lKOeg1KjNFCw3COkb1CmoubMCp+hzYtPYuep5Haj1SvYveJBLIvh
3NMuS0K6C9VwjCLwjN1gsdZO8CVgFdyPFBi9lr+NVeWv1Fq0UJSnyE2ro3eRdHNzHxjv2VK0o83y
pGUnvhbXjNUVR45Ee6IHXpcgOF2h8XMsL7TPNHFnmYu5Q4KE2AsA3pj9Lw0JU6sIAMu3qZbfLxTK
FNY1lWmoCE85l3nSAXhJ3rN3HZ9I4CF/ytrnHMN/SrPVSkHF1rqHohDd3L3LSOeYSNIvkJGo6KNn
K8GASvThbaTUU7A0/itXGtePhdxHkUOaQ9aCjTXd0F33Zj8NOQjK/vgwghMJEQjB3VI04NcvDJcT
FVq2XujzUSWRWppPIspHL4x2XGxXCW5Cm1NURM5G5vLR1COSrlw8LDVRyjVOa7vQ2YjFnXi9teKr
bzgo0mvPLrZYaHHfcaJQCg66TC0D39dNzYaxL4UqGclmejfKk3gYySJ3E6eder9b4R2yhOEx9AHQ
+z7RBdLqPYTx04oASl5a8x8kPTCJmxfJtGr9Rwx+8/1t9q0f1dNvIonUufqT081V1gTVN8ualWvj
DwAOQ6oFbHENhBQ3/Os+nGzj1tc+HwzbFbN6Wmy24JIR8Oi8qSYUKyjoJ1SBuEoU4JM8YlgLE1/v
b1ZBQeRV9hEXG1fTcSwH+ND2qetY8BpgVyLivMF/8pLQr1LegwtAgrKPziAXU3eYpLfJPE84/k8E
wuPO0nb6TB0kP1aUktIQJhG8kH7Il7fRgujoIGP/ZfGPizv23S3Mnh4MVR6FnUiubxFYKaaqSISw
tRAzPFiVqA5Gb4dbNvPrBZWUJUAZhn0EAFn6eAbxetHhRnyg+tV9HguBOaDbpvdOMSqciaWyb/E6
DTTPLJtxMxSVtNYFLa99Fw+4z9vgvfDrSNpPTl2bjd6ZYT48gnHjGo9nTx66uFYijfeoZNUOQ8uU
mf8KI1luXBnt22DYt6CN8r1aLhVsFMtBqpp98QzpS4ECFnmOF/aqcITLHT/YhN8xcSjAizqvVfys
0hfjhjqacCGcgV5g/I5oThBWfuepMyu5yumzrkhlCpjwtkGywRnCZDj/vEOCgPqzAETeW8Mk05Mz
41fgb9J4uQkBuOANi5/uq1iiIbz9NC34zaYqR1Bskrb85d4Iik5eIy5lNk6oPx8vqUUe8XQVeKrM
bhK1ypAYjRXPduC4NYkMGkRv2V7m2GdXcP9z+TQTUqD1z3AcDUzmJP6ZdL9dnifwcSafM6YNwi4v
uNdLx+BWFln3aM5wK7OIFc8McAWRnpCMmbFYi4k76OyAZxMVqgm9yt0Qf8m7f/PA1INNnZ5LnXdc
868CyGXLhfkJXj/RthuAVIqlWX3docaa3ym9ZeiIb7UqZIMPht4Cb6t8vCh0A7BwarHSX04Xe8SR
ItjEVmv0bskrSqPIVugmh3R71YJmT+ocXTZjpQgZVZJH5VCif0PV8WhUAV3qzOX6+7zxDgOdyYG8
9FsB7VhmDBoy61cwChk0DdQ+5++WJwlvBzn9mYqBVMDV1C8svqYJ4ka1T6+99YnvaTEX5r9vmKtY
7tF7tC98W7TqRJhRaC/JuuyPPT+OAGrg1Jyt7ZSQSp4lyUJHI1S6XzCmDzUIEh5/z6qHk3k47dHw
DNZOK9tCerCahPSXkFPDd3W8cUfJzY0QqyM/1cY+tB8hkbTy09QL5aAiUWG5buJKjwDWGTDck57G
frJupQkIcs8Ngyk6HfZOjPeO6ej/5J/Va4Oud4r5r74VXYQre4NsuvSx1yqbBu1nnE6QnPY9U6Dk
lfQnBx2kR60aoC/B/X3X4pu6F2i/8X/pF/Q7u5ShLSYFUNn/gpHh1qZVkwk1igHX8u4bvVRV/erM
/nkA5N0QuBz1kWxu/9pj0N59Y1+nQsAVcwZJqlR4BEA1nWRkF4+uape0BVCUmokO3ZDk+ITg16c1
AF6CRuk5kTLzzDs0hk90HO+KDt0OQQPYhovic+kflD+AjO+BUbS9TQadsXgt/z5Ewrz3f6QpHFbs
tWCcdI2jqT1eVMDWVrjREIuxYS1UeatYek9eM0gnQ9SOlozqULmHfIiCrMtOyirjsnURllJ2wgPt
cPfzc1XYaRDLOQOc5UsJrDt+FLpRNJiOS1v/Q7oCcziQQB/wA/HUw9tHjY0hCnNmx2g5k12DYBuF
qfUQ2/me5Yi/jI1bPXmA6EplDy8KyLQgW4WyBSnK6BI6oKVIMPSUt+FJPEth6DC+iUIgqVB8AwOj
3uQKs5MvG26RoKTbiCAz8EUew5deQlqEerk93uS8F1xoeteJPiTNmwOH9VsDSCpCoF8zK/Hdsej3
qPP/IEJh95FGRiPos9Q9IRZiZRwVjzP4Id/FjkuYW/jsYQK+D69ZDU0keP2iBZV5tMMV2u0XE1N2
j55O05t0cz55JdqIG6G8XxOuEQJD/sevuEuax6U6p5Qo4cWr81MrZVUjzsh46POlFuYtxxkgPJhS
YBRyq+2e7Vd7pXqYvFInq6ydSdcmkReM1hz3SPDQNTiWYSi8e8+c88zZLU1E3ZGCUsko4Acd8oes
kf3wYjbtoYkQeBmStNJI77d6wYrED2qV+qDMMBFK57YpuYALe0qefuydBtK7k5ysLow1wLcWXbZd
Qwt94VtxNC/vw1avjr0Fk/YwiZG102d4DVFNzUi/HB/3hasmA/FSBZea62DaA1HLwNZH9kTMhM0W
XPaOlN5mLUdFtgwnUI00Q/SNnqqZhC9Qony1+h3XAFWitGSSnyBlumy8VgXQbNmMadUcY6zIxKzT
BDKajJhUBZN3xf+XBGN6cwMdnWtWf5uzbCzrLynXN0Vv1MSnaeadZpcQSneQPB1ksTbeF/r6Isz9
xSmVIokaJedpSfAEcFAI6lL/px1leva0jUUOLvhJD2s57p5Xx4YB2Vj1hF6lmwyxlN8hIow8g4hg
SscwW7IiSGor5/9smv5SuiVlxaJiHldPM0/UTo3Ng33gDGpH4SG6MDqDYsrgoVQEns0Af2AFECGm
8OkAP78M0eHtnN0lyZDhlvVQbPH/xVULZx0IC2EDxqWRT6RzqjbedH1RjTptvVjO9CM0vqWeLYi8
6Jq3D8vorH70pOC2lod6qqCMZNl9AYK09CTOH0Uhdb0um08tFh4vBrdvXl0ERWdJ1a2kQYTKqY0r
ZJCJgZMBSwqLccrBzXJAIOejxsiy99uosOi+km0GeuDZdhcnv6Yz7Q9ijybtLMoDmSDcgNubXavZ
QJCmuJqvdm+m9R1WDQ2q/Pq1QUhs/35kQTWjIcnnUvOurM28evR1h9rygWlHEWIuXyUFVe+MYsi8
3G3/ovfAkkEYrfg5b/Vheilw9ErMMhmzoFSoiba0BaFpL4knCYR2PC7r5hwRHhBCCf6KiGrJrzyU
buH42A/YTqgPk45usVhzEF/ue6iKO8Dcerm8wOMhop85uANR8Hkwj9zY+JuSsqSsyopZN8gHVV7T
v6wankc1ES18xLBv1mUokj/j/jAgHwqB9C8Sqd9ovhU8nmmpKtqzN15dKpp4OorZ+CHCTL3urg5G
t0yfaGkNUjFTDWntEliYoT/aKc+xEv94UZZ86NZYbTC3mOznQtwLDRJ2BllafDWecu6CWokts3el
THzG3uVmpJwL3ESq8PxHQLAY8hld0BFGVMecsk8RZocDGJDinC5snUW7iYVz0TvihCWZEMeIR4KY
KroPu1pgvRhGKY5b40nLOOCTetIG/0XCbZhkjQ0tq0hrO2T78ABwlmnKgaF3jebYZS5rHHifWejV
kWMHhIGfQinsVXlnHVra6nDgay/+oKielFgZXclEyW+LSoGOgOh3GOLRvctTIKuV2wHiamrtfzhe
kJ+nZzHUWPO6Xz3bIL1IKi+Av0BiFTSV+UWCZiut/okr5VqQzYx8vs5zjK7W0PfotRYe0JOTFokg
pD/YwMgPp2eQtFxU+/bXjfZGGB8l8ElMB/LBGe9QcB+9LspsYscL4V5S+lNNUxab7MmqhtqOY5UE
DmOJcEZMVPZ3S6LHPzUg6hzksh3Neq6H/TK3qR2m/uHD56//R0JUgJdtir9zC5k7Lr82aHaUGwwD
PVppw5unRpTAYAYHkcDILFLN3X33JhhDS6JexXvWhf3bjX2KkICKRYNHRGfabVRkU8t/wrezJO5+
51B4hoLcWsFod2BCWJcZO9AoHx6QE9wYWmCcq7uwBiPzd/AAHRZVwBn+F7RrFR3goYSKxmMG+cl/
LB1WgWL5rQL1ggAlio1aVgxm6CHV9mS08v6Zvq67zNYHnRN+FfaeLGnMv7Ryy7mgFArpn4tiLIis
MYapFbMUuxN5uyd3W9PwiBSIEzD3fR0+gqAFpCbFVL3JA/MzwCe0LHP9mu4Rm1D8pnbZTwrlrXxQ
pdeNJEyyvquTtyh7GPBZz/RA/65HQtdHULe6qo9hkMEZZ29AdFHV2H0wgW1pQ8y1IGguxRv0hFjh
+Xqu0QPRVggXK2HOq88PIN6yIf8B12jSUImt0lCOCAK1EeiDSaym5IMcL5Wo2uDcOQO8b1wuH8nB
FG2LVezaNreWojMhwoGKokm0w9VYv2j72xaEFPcjT3NBHj030yaYnfPVIbjb1kVk5RsRkkCy0jTw
ZgTq+AGg8VncxoVN0mdIWUnAGQHZLuWokwPJ7HCe/5Mkfjl853KzELxSk4qsvMlO1vMtjGo0V2uA
TFd9+XEJsVXo0KDNTAmRQWBN4rm8cPEyyPBA6C/SDJBm7LF3JoGu8FQxLlj4xAZ7x7iSxyoIU0oZ
CyUlM6BkZ7RMrr/p8HX9hFceX7m/Q8LUXyZjyTBQxm017yNFUf211jOOxg1juANO362REr+u9V+9
FjLP8EV+Rm6kKWLzPLLSvJjILVs8xOI+sZZ7nzaixURI2tNlQGyHXrqSW82Dib7X1TSCupqvvMWf
W476CUeuW5rdMxXjDXwoLiL8Q+ZHqC5KJhZZW7qhPIpTgg7nz/sS47h030sYZ5pv1Gj3KvmC65ro
FVSFGTlGChmM7/6qmMFG1/R+7bbPbFjE+it421KvAouueXG6BCSLXlYrbHYiZ5RcATJfCY/9bXos
tAUXCXsAzz4PM7DzjBCxmk/ihMEFUYPBZcujlOn7GfyTlKb3090gIVTp2Zg2Oa2DlTsgUgPQK+Zt
BxxGuMHVlXJlzETqyfCOnRSF0vuLd3HMoCQUMOlhahAR1cvpeSiKY/va0t1boKl6ECASomWxPBVd
oze4iac6HkxchkgNx7Xfwwj7GZmUMVqATxhLqK6pwlVu98Xq9tXTZ73vG3ykoOB4dOWQELW6nM9T
dpV4s4sbdgzO4gB+poLjeAQl6XCVxFR4uAunv8dPPVnZF47oH3lBJUzB3Oczvzz+hZMaK/AK/VtB
tMniVNPyt3QERBf0EgaAB4rrxcnzvaWqAzTnahdOqsz+dfBZ7jsjImb1Z0RafgpF/lZX6ty03Xub
JOYVyLzMIqi1/HzOqoDsXQPQ2rUCQsiq2s983NJ9OdgSIXv8ETn1C8uwmiHM6CnbFUBDZdqb3ALm
dkH8xu/Qhx+KtmcG+G0yTR/ci0mT7RGaymqvaH9tkhVh0osbknkduT8pnuCiJrMmleaDOI21l7lC
7WCMaz+/0radtuyJAM8j+hVaozmrLnn3D54/JoqdLWfV1VCHZXePBZnelKsWcqz34Gvz7Z0t1J9a
2cojIc0/go19XL8/nWtzROXyqniSTlh39HdWowigyHqBgWmEkCclS/Y5rmggDyEK8wWvv/hM2fN/
KYCgxvQ6Zs8VHkAbRG0ETSEU7kylNw/2tCy6mZaYtBnvRBqqhMf7Gk3arGksRtDANGRd5Fx6S0va
y+EBoKARNIsAF/N+1qgNxFmRWBuTKqjVnLysHw9IEh2cQIR2pqQ5EGhMh3kc1sid1jAi0tAQAbXi
Exu8tlRb0aypL5Y5QIpHmdBfHHyB4YWkgaMKyzeXRvs8GZDIg8o/K+dVrQNDSxq4xVZZXT63RkCF
Zpl9o3+KvX+KBN1Mw76yFedf2w+leHhunW8ZOHYYm1LV1u4nmrd3s3JVqxs8Jq0Lr8WBXSWmRgnv
QlCplqwTfkjcRMyhriX+jPSgX1aJHiiuuorTmUE6dvFPV/u3F161p6fIbYq2YvPDL6/3TVfl03rh
TE3Q2mRjoo2y8Dn4cscjVIZnNQof71PwxJyO8roGG+a8qBkGrX2xCz52wZchXKfh93CJ6SlXCg6y
v0G0bf0Evu75WzYoI/CGUSPVaRMyUwkzmQKjg0RrWF2SLkRLs/C56lRwtZrs9iLhTrkva1Sct6lb
mBQ7NkGzSpb//M7fpz0NBZawjDzLf8fiHyDABBSrn6SoEEUe7p277oAKBIot52RSRrqQHg3GZkJ8
1oODOKuvmh0GE4lcqjN5uTaKpssiScCDyMLSaCQV/pSj8ZXvPUQIJzaRe2tX8wZb/w2b2vURiDCL
X6wxg9qEvkFBZnT8xYdoc29kg3Llzo6gKm3r8z2mOEm3jt68frl9i+qE0Dn7avGUfLedV3pkSHf2
7GTl3VYlou2//wl/W1ngYX6nPXRda1BYtLC4GC24vklRGA0vGylWbxUxqZWb6HIOT292YkAqcIvd
fwmFphSxZcaqEeqz2pRViY7JLI8+KeRo4ZJHCjsKe6QCE0aD3aVenPRNOKd1Dy78scVo2Vu7xPjo
Aeql9/vQw0oDnGQoIcqWpMoXZh3eJMwhQRCWwWYilSb+NF44Iv+sRX5NRzpcjFfDV3D0g/ZTWXVj
3kkvIWbXlgr8qWDoPX+DFNm+CuWowmmkUKUjFN4iT6zTguC3r2wjDi1oH4wlYIv9GwzlhVPgWQDR
FkGGOtk5e7zKk+UpTf2mUFM35TEj9qAFpPUNc9wOONbsKp4UO1hmNfwXlaHJ9fKOQ8NNqVVcS9Pv
HxFhJ/5+uYdwtPdmrliRHPRHBZ5boHjxMilTWDVgZIXLEqfabLFrIq6smkjSpe2L5ydVFAeY9+xJ
F0naisjQekrJUhiumQ4whTmCFXRvx2HDmMA/N/7kDZciKkuIPLYwnBYOogrdCmO3ybUV5GtOhdDI
h7BNHbo1Ju/zbU1fwjHOI+lu3su/0OKQQsCxqM8sUdtw7bWLfflJesgk3NhOPPugR+tgCwmkz5zV
jzdGH1cUb4DFhsQLWPAcNgFMdDM4V7yVLSJJs1KG3IGAOro7T5L3VL/fGHdONNfN6rVXkiRp6Nl2
Bh1m16W61ntlUvCxgXT0MeSbHWkBO86U/F24NOgHFd0bwG76+jIVmeEc4bWe7ly4EUFgunWjCn02
mi4AqxSgc4NvKsq+v0zJp2aSbmdC7qla2qmMruu2UGTFq7fS61Y2SvRRnsTUwEWPDwSuPzMxdDvV
vRy/vG1JkAlE6RP7xenezA5trmPqiMmnRzemGRTo9IOD6VED323PRffp78Y+PEklvBgmTDtXXDtK
iP/3Bu0U0uiv0m3641G3lcn9sZc4BnwcFSsqoYHocWDdixFQHj2LXqqJx8g4ZGiZgGCoEogRFrpf
MKDLAuuNyKyJWUeD7VH+v5i+Dbb/hOX+3UG/hUWr/PqwreQ0BzhnFANMFFO68EfbEr21f4r5fEuq
N9h9l56bD7CjNQdUUbnSROy9lsBqDfeTzhu5QN9LtekDZljFSJh/+bX1Ms03nvirHTBG5iyz6N+3
3n27qm7uLODdX+H0Ar/MXP8HI3ul1cD9+an/uEgGh5F9uBFpcTXing2iNfcA1lPxjjqv201ZOA0a
dq6yEJMhDFnQ5yk2OuSmwem0RTHS3HK9eIyKIFuGdgFhAwCPNFNWnHHiWXrQvrluje+Cip5qiprx
iAUIlAnrDHYqGUJ33LiWpgrh19V5ya6eCKu43pLohFSyi6fbeB+zDvipBFWAbrJBYZ5xce+JLYSl
cOproOuC6Fc6zMnjeLpaP6gW9gq6+E4PAsxj0nuBkmAPtoIFesUXAoebkhpa1ngYaHeHqwvr5647
Yqvb1oUipkpfISYs9mBkVSLAMPHBdJ1OdfmXc2Sx8LIMVO0rBZELVrMp1mAEiEhB8c9J2hWqv6Fe
2iJGaDTZso0u1rrr+Ib03QLiJmNh2Uv8rba9ZW+XrXbC1WydxnrYABAOcjxYcURI+RRXGF0TeKR1
6hwJse7YUJ4RoCflL/jYJOFV37ztFZObvaZl9OSAQvnFOmIUx+kUUJCVJ4rX/CXCDTkLZezSTh/M
GeDcbOgms3C1XazM6duafuHQSzjeAf2G34P0HDbpLOUOqwuhddwNcRhaq36NDicLY0gFhIDJpDcD
73LWsagNq3KD3vJ7Odc92U4fONgs38WJrOobBGeeysNP3S7+PKcut2bJ+I28zDaLNSwwNAOp+FM7
oAADxER3/sEPQyUKvtLAqvDLxrULFca2XWZ9XF8WFdysPXh+M23YTgYME51EqZTWd2J0zrxaQL+2
ACcC8JOF+hTlBqp5T7RN5ufvje5UgVPM5kKji7kxrjMBm8kLe6PiNR+FT9Bu9IR2S3Xz1QVQYBDH
ERQIBksCo9k8vaAD8pST0ng2oM+89XnbsdKJItwCkmwVutioWsz21CJcNNNlQZaJJSuOCHPJayTf
+kGmIye/7MmiPF7t+/3VTsx666UZJBO9T5eSy7X3cfiV/0wgrtMMN5B988BaUXExq05q6eEC5Kub
BscjU0nFGImsTd7CooaFioIpyMN2tzv7XyYlhYwzPAoVwJC4dOLD9v53u4Ye1fg7ocgyb/qkQkCY
m3igEdnHtgNUqQ4cw0HdoKEXfgHdkfQ9NjGG40+ZSuD77OeGDgUsrXiyDUXLKNUOCZXcyw9BhNHS
SvItnZjYoEH6ztPvkzoIgyUwWyAsWYhJwlTIYcI7bPCONzcpMnjufwpt1ougBnKp4/1nRLEy1Ah9
egiszxCcQFGUU/9cw7QVXOI2VaTZL2haxlUQIj2lRqmtJ3mzBNKqmYUtdR9zYNrh0BIWQukeukpq
1vFb6hy9iwhst3gZXDzSYvI4CrJGPdReSAUrVdnYiFQGatJeEtZilV6D9gBQ1TMykOERsqGTbVWK
iHDtwxmiLc1GVSv3FW6hzs58wDlNRZUXXRyHfY3TDkXkOzFxE3ZTmCAGbSfN0xOBTCuPj/pr4KrQ
GYwTpD4oKmcWyUwyaO1pU9sisnF/4pkBlHZ/ZOYlolNv/WIqG54/1dp/T7J3yAVjNH+vCfl81EIl
5kxb6Jv6J+SKtO/Lb8bvjwKlHH1GzY8eYvaVgiYu31WcY0phXpqQIuikoPg+nECELhTdyQVMRbN7
XR6qykIOWZZHqhPihKY0dB9Ft/4iA4pHcETyWuoDkPpCz0geh2yScMZwQfWDEduXXfRiFGlKbzmA
vJ22MMXFtkd9q0yQb6pZN3gbGaHH3WEncD8+qz9vpI4uQdR1JhfqfDqv4cpMx3lu6e2ITfkWEsq5
qmzC0g0I+OVeR1lo8la1gXEyUOqfkgLfIl2CpfG/lFzH7ouLbkpupwZwsh8o2bDQNvlE4kCxHplR
FWBFatysVabIIdpiG3UYRxCRqIy131CRKI9X49+NHdXBbgcM23TNJpP+EsNZMZgVXr0nHlnyH0aa
l31P+ojTbbUB2UsgByVXoZpZzuN4xJHYGd5d2pSdzLmc/rU9u0LhC+YLtHeAZOkx56b3P57VR3nG
dxYWfBmoV0iUu5NprHl4W1cPcKi0ULaGChsF6sNgclyCYFXq50CmON0XT56P7r/D8JZ8qLxAwAhX
sVmBHQ1T4b+3VhayTKeaz5Wq0s2j466To6Li+Xu0cQVMxU6XHO8xiwHZGaBHtc8P/AwUXnY0923a
+p5BBWsuBvt2DuD725JmzkK3iQ5FzBJ3NVXeLcXv4JqQd+SIyGlhhxbV7PIrkLDdJIaoqGvGNCN6
e8FXP8P7mbLLh0MGkWb8+Jbcyfax5I+hT3aZG9qUSGt7UP2BOvlXsmqPb02on41HckvVIpNd8D39
CqJaJ4S7TrwsSBuL4DRPC50J2E2pjxtoHHCURHrQxEI/IFkI+yTTfXWAEqfQ+ftnX07z5fYYplIj
rVtjDGliJFDJjB2/x/b7RJ0oYRDNuwDw/2HipwKGHGXR5DKkU6eYYJJRgbl3Q6jhdg8mHdCdZX2Q
opQGqbRO4Ak5dWiULgDE0M+DLKxpjzxfhXpavv3GcG8MKY9z4mxynZFDVjEsH5pexR0R131CvR1b
DIUiPmGJWlCj/swnL/EB8KnMdkkDOs9CJOL2yhUCtg91csiIrkxR3Rxs68sRJfLuqyyhP3dRlQYQ
cm2PRwKykfyAF7OQJjEylYf5aAegrSpitpFzMsQEhhntx8K7Xxgjoc4wII5LTNCNmggVHZ+YRW7H
MgN9V+aWJrx8A254uxd3VuTklNNy/5W6eaRlPg8sAbpv86fd/fCs2uaQYtHKDQjyqVt4PBJz9hvT
5ozb48wRW5Xq4W0y20h+VF4vb/XZ6ok/AS3ziSel020QbHbqsYaaSMy+hYKRdWsFL9JvqK+G74xb
OW2HZcHu/7+U6eDSAMkajira6JW7cWlSEwoTYCLsgNBgMa4tJPaJn4tL2ZRS+9UEuvK4iuWBaSaW
lIbf3ADZ+d12dL0POSublRg//0Y5geES94OGz+OV4bBHz/lQeMRLTU3NdGiYZZdXhP7SCe4eetej
6RWMtBepI92zPzwumKK8T/PYi8HeRn0Ml7MCWu4+GoBl65++gH63hezTtu8fEVGyWbltn0cUJck6
Y+QDbMmGWxII0QmOAT2BxkrdRBZe0GGgX87hyAw2F5v+TG2VRVsasebe46Ng6/tRjgOlAu+gqVf5
EaEJVb269cLFAQ0KKx0wjPRVfBVoqj2ydQkpa1Ws2bIETO01T70SMGPg8XVfzTQKy6+J66IxV2dz
PP1U3xoMTKxj61Ml73i0x4zxn0YlGTjfnL6RrkgjZ4K+DKMpoWBz+bNbGRl4QxYdvvIXS4WMasF5
Tgjzj7N2XpoTVuf03BaioeVZakbJKEY3YLGxOrx++xrBzv/FmmQwcs/2LFHY+0EIL8Fv0yejMDSj
pG4xHTYAK3kfQWbmkB3QXZMqlLzgGVapLcgkFUxRZtbYUi+Ib68ON49PkOY8zKRiUY01Hw5uLA11
pq7xv5vShzLqo50GqlYQAY+aT1Is/pIcxkEIKB5lZWcFXut6NUgDoU+7DDe43G1zbKKDr5NzHBPi
iJuSC7X+f6LL5kkREkxeRtK1lT2161SBMydF3h4VaMDHE093GTwS0swxMR/rkJjXbjoxjo3RaWOA
WQyjgS+vZSq+6mtfBnyFydyfmqmud5ZIjUpn1phj1nzJqI8eRAOVmNuQogU9uLuGB/YkW6CT847G
7kRllTDHNyryue08DczPVzeRy2LWpoopbVIH7+RTWZvXpnHkw6so0SMhVxtULOE4XaV4UsDkcw/5
yyK/MhwIthMVytJei01L/1T4QbhwP3XRnuE546OX7y1Sj5eOW7293X6UtKGQphPHQAt3Kaca/kw7
HaUAR4lqG6H5bOvtVDMJY01Rkyi59AtMFxoHpE1963fyUX7/IcWldcrmxW3gKdFynCWp9rVWVBq+
iM2L3+CRTbfqeQCMH78xrJCR5Em1jCGopO18u0XM2G+js2m/VIrzkV7QdqkMNIb6ijNEZlNtlv+6
9vxLd4MTPGZ51ZvTo1l4HYi/Jb9uqH/I+NTqIRkbWK3KksHwuyVgQqVOrvpHQqb2LAs07vUzLyL8
Gxy0UjBGTMkvfJKOnK3Fdx3fhei5HWjm/JLxdTZ+KtqPj/juVAlHs304Ettu2hlwJEJTE7Ow2cGv
Aaw3ouu6wQFkieYHc7C4N8x9xs7+d/YxRZNuF8jtMsV67j/rZD75XBAYuh7eFjIUHytwmA3xg1lr
wpIssuPqhCKKRqmSx17UEFH1YrlfruK/Q3n/HlyyIfuW8tyLJqJQ7DbvAeSVfWuUwwus7mahSd3G
m3AjyzBydyfRdjsNA1TzqOUT8ye6oc1XeJTzk1kZp1TVJ3EbwngHFhTYV7xhQMggwMIL3E+LJw01
ss6q4QuOJ/KLpSU2hQxG6kmLOtDBw4h3gr0j0DLAFVj1YW2r3uKopZWVywApnjhxGUYoRs8WMMaM
L2B7kUw86XsGsCxrRJhdr8PZ0cz16bYgdF0iIYOfKsMYw8a0cHJ2drzKFEojSMLGpNi+mXqjBTsZ
+oKvIygSrOWsa41zYYQ8Df/e6sm57qd+THECUD8J7goDsAeA5hXKqkd6N6F0G68Gmv3BgdXMqT8W
HZ/nWVTSfRPIsXKMV9P9ZPTZ52pxnBIz2ELrFmoZjHhvGRt+Cpw2t916To6upg8F/0kfVicnOL6w
JuZCyKMfqXqT4p880p3auqDPhpN+U/Fefd497yCMTsLNcqrQmyS/DqUzg+k0ksEBL1luU6eaJUlA
KE8CpGdakrbI2CF2Eu0Cj/UbCB9dJXYzeg6daCToRp1RXHcjjA7KRSlsfSwvpJy9HnsrNrxXYKVK
1U52AVBqxALXbD4rAm4HAZ9S53INd4uuPGajDReAnoLPMMzfj7ueTqP4Ds+4RzMT5D0Em41p2SPE
wS/rgWKxFv37b96+ymm/KSQdYbSL9qN06Wc2r5WMoy9KwLtk/Zp3nMtaV7AatRUFuOOHlE8jUkI7
5Ylsk4VdZTgNoVBOOYbNiTkDDvRKZ3qkD4sxjqtrLjYGNUAZqNFosjDHGvUuAb5A2mnXxIXTFs39
S8HMzkyx3We0D0Cqmu2L0OrKQUSiNafYB5FZknS/T/+gSeu0uDNNJeRpXM4cwpmgFpnBUyibyQBz
Z6y/Ghbxp+owVDTRGgYM+lAa6dmPiAzwbqZqPLXampyNSgVkecELaYpbyJ3nS/dS/iFjjlZd8g/3
RIBqOI9J8qIUBR1cCpquZlj0Hl7PcOAMw+HTN9gCiCVfn1/i5qtB49mf5an211N03N3g/m8rvDTM
fZXVuardrDiT1UKdif9idcND/GJ31pvcreviZCdrNfxvMxBTI9WaoMXtR6wvz/ENZFNsseXHsH55
35Ksy4jS0mcaX0pVxj1yKqbngc6Y4FQyfWyb97OEDkDMSgn3r02wn2RXOjRaZeyR2JJm+kO7cws1
XbHF4Am+FVPqRD+MQy845VpBAu0RNA9W83EfrwGS2ajbO7Du/OCgXL+H3bXJ0D2DHatG5Fj43EO/
BUPUGqgK+JXQDsmLfGe48n80fqbvN6OEWNTTRnP4il1/a33taZatUpHBH2d3953QnCj504ZGLYvS
ukD4VtN/5tJRakEBarSi7YC2ZLef6RD5eGB/OFlXzi2rmaGc/eNFOWxv9j6LQLrPzC3v7W/aoXfA
Q7dbHMLJN800TTBV/Xm46WBru+/mQQy159cIbNpxNuAfMxuDUhU1txcq8gWK2+ksNu4/P7pVJQ7J
HQcbqs58yFR6ePYytnQx4pnzeQN5lk+3rmUPZQNiOHDMokXI/yfldrzkgUJfWtNMNYDA4SUJMqce
OXynNGgXzeh4Nr++Bkm+vYlkcZGKUJEGW/cyMW52EUe/gTATLfihw3VXJEVQ0tu61/V1YCBezwJZ
xm9sWT1adTiTvHXZwI56CfqaE77XsfpFghDlQ6pfRa0gK/m4mBCO2pleW4gwa3d3N1UIpuxfNOiY
XvKOHiGOiyithZh5ku3QYvgXEE1doUg4Zw6KakucNnFzuA7r6VRUv/NWHGPO6Q62L24SqKe6jT0U
21rM8mXN0E3JW5p0hkjFACDAPEGyVBLZjhpPh58PCOiu7wxqPi36UOG7bx/hJ6BhWGahe/PknafR
t5u1937pAh1eE1ZHrWHZ75zP9F7Xaym39G22qEG7wV72Zy9vLEeQuWGWGBqgjt1mhrvvGYA4YWGq
zgUJ9HyLuNkUxY9gCIOvsclv3CIla3D96wvqHIuZ8r3WNrUD5ZWG+5yanU6pBlvJjv98IAqYBXY4
caoMO6VkYJdZGVJjWIfRHu868YYT9WSxRRM7VDMiN3gptSjBQ8fb+DDdoPCtwP46I4MPutKxn5w/
J1NuFp0eqndx9Rvswq3e5aL1daaxySMQM8os8FNPA0CXK/uvqygZ0aQ+Lp49aRwcjJ1FbtOsNE3+
Uce9UwtNpArc/at+o53lOPc/KuZGrxhnIP6JHLmvG6ytlEqvBfQVKeRBUi9wTDtptFm94dzR07i8
VR1rD6WdOg2lJROITNr03ZEoY/qFZZe5t1hay0hPoaxKOul3WW59SE5IQHwWUiEog0zf6kPp9tlY
t0ns8MUSdYwGTr8j5FFFeBHpkkANtBhHucgxDaB+bG4Ci8+9WnxnMJ4MLzpJpD7yjgY+tzncyJi0
KiAJQu+fW9IStpTUILmbJAWT5tAa2MmbuI6L8hLWKLt/4CvFcfoboFNXqu/9XAbUdAWBQ0T53k6k
SxB8h0hIEXH2kmt0Y2ApYGxJPXSVbXlrCr2e5c3aknSg/Wo29FI9MoTrerwv2/O+jVvzRVwlYsyc
atGBWdXex2fb4uiS/0HDDuE/dh9LqE7L2RtxcouuIe9niYnMyOELyZ6Mm8xyLIP72me+c97ibabS
NbO2lTUNziPXtY8Fr1AXcFT19anFq6y89Sp/CmKsYcqgpw0SONCI1Lx7GxMVu/1QhIOoJkFnDq9s
3079h9IpaC9mNGh+lTrU1112wkH8TZp/8Wg/Qr9ruYFeGt/YD5WD0NaNtjBQYOrMnvgGZqzomjnK
2t8t2XQ15jLo6q1w3cn1CI6xW84FNrKRZoZsQNnYbRRSjTimWoXSwrVIuNJet+Cl9tc7IBSI+Z0P
OalvAqks9tJsD1oIOWyI/JEnfOPuVUijZAa6rSWcdqRe9cgHJf4truol+eNT2an6pJhNMXitASU5
QA0Gnr/s8QcEQ/XfovMlh/UwVBFSVaBPR9lCxT4NFTpYvWfJT1t7ToqY1SKvEPqmC09gQuLN4Ke7
Mmymn4pWVF3GAtQcBmQQHk3VE5svfzIZcdtec7bxJ58YON39Q75Hh31WPA23q6i+ThcBrtcHjJ3J
kdmyaRpfCpD66FzZyQuBdfeHApAIN+yiLNWNbql612e6U0vyg3uXy8o6OqgoB5mLjRkf7mFpi43Q
Yzm8j7lhOVnzKZf6aV04ViZf0Rxo/dOK4ko4eI2xHcGKRj1L1RlDl2ExPuSZ+OvZHJmsBIvzQcF/
gseS3dHYsFrh41VtbGLbJrwQn30OCff5EbNfl8EGmgniaAEbe0RvpxmU77JBT9J4z2IV0/4zlbC9
5UI9Yo1NjEj+DPpm10cGjlw5VpD9wL/iYW4k59vTHSGy/SZ6Z+tXsdC/4wyEGXQoZBonHIFrNL+j
ZX+JyUVdhJmSpj7xCfAmYFfPb/vscSEX82RzW8nKHq01dV8jiHIGw9CjtdIFj/Kq9i20Ei9/5b3I
xFJiNH4aKYYrrBlO95iEVYeUrYqzG75CC/bipYPcymArSPzhA7sCeA2vi7I7CzlqFjdWyiTjX5rg
wDGm2r07nnATf/K45jxa1AublOo0FsbSTxdhcCSWhTHAX8s67GVJEanIeyBEZ0zzghnsaC7MM/rQ
KUEMIT0anzALBGumPRo/qkWW3iq/+G08Rp8RU2oIJfe8e1kBPJYpfZctMxBLHaU0C/U6b1z9d+5h
AxzyGEAvfCWfeUvZ+QnqVv6+ezPxmqLzRaVStNk+NetXMSo8W70e1uzA0gZB8DnaKtErBivV1WlK
99snc+8XZgD5YmAhwa8FB+fSzfdtFG2YmxLevoInY5A6NtEHfDt5jnlrfTmk4SKbSHp2ydUHsY1e
NaLjoey4kpRwUGWirE0bEuTqqCCQ7cPFzVHIz2m9q9Z4NTSp2G9cqqGhexcnOU38NMFsEq6T7pt+
HjNVJr4IFpCUybHnkSOH1ZCuMB704JdUWUN0NII/QRj2X5H+kTOSFRetSTT2ToQRpt0tuhjvd+3F
cd0Zuzcc/8uamuYL6gjJIRJmFbBUKuy3qhrScjmD7CydSY6tWep6ib/2yvqKXxKL7Zo0U4lQSkp7
5JTq7IAG10gYmQgmJ7T1KX0CC/6JHCcw3Bq3KkTEmVZ/PCVtb/bHkabD52EkvwyGcWmCWIMoph2l
NP4K26v9kTEV/sv/lS2CMabJL5fZTDDayhn0t9FdcaSWCpTdKy9gShE0Ww/W5DO3S5UTBaD7RodP
fclLUUSo7aA9yO8GjXc1t/53A/Z1c+s4dh7qa6sHsZQwXl/ZaMx4i8xoTP30V2+UuNAbY8w2y2k6
7qrqsTzZfbKNF/83jmhcYNLSPGAjyuKG/MhCRa2oH8IKPHw4QRhDcE7oY5rd/labxqxrSyk661Tn
P6Pn5zPnreuYaOWBl4sc516dCvxtGqeqXLHIfeziwXHdAQhWhNmJOmAlpT3TjTaldHmwFSEUMCRF
ALddMfR58EWWj0a4S/b6vZDzjgvCiZ1osPMB72AoccNsZ9Ftoin3NvfVQRATNACMmXXW2rc/TCuo
waS6m+0x1O69zXchDZwxLnnkw1XsoPqXjgBz9jDjPKZnRLIAFk0KuhNw78SIwendlNVWd8R23udi
7Gzb2m5PQbfjsLUX4c88rvojE4KcuNgLw68g6hzV8/V/eczMoF1WEaig590SGBQ778xaHOMAhiNr
vbX+idKfit4TGcQC0MAhyIl8pYZd6qbO75AxbR5/429b8WNi0DM1H94wp0PsyDpHzNdqCA/dFff7
X24UioPQWLQyknzo4E4efTJl+1WJATNyojX8FInqdJ8ZF+UvqCdpAjUB1Kay9B7Of60KE+FlCuP8
vxsqp0YWgeCTAy2gxmUAQoipdlB/X2lK6+ccYc0sXszSai+ReHZSaqtY51DCJjiISzq8x0tAe9Hq
64IPb8qEWn1jJj+1kkJoMhP6EqYDVijkopVJoYqu/bB+HMAMXA8pE8NDJ11uQ7KBEZeRXwGW+d8o
dYe6AHtO5qFiiKsIxBJvOwdYQCIlXtiQIevX674VFra/BmMU43Kpe+l0CXZp64t/Txph0JW1wOSW
ipSSbbyzDqNrW/Oclwj1QmhuBZ9s6K5fpCUdh2SAkfLsodK+UoDrCfDs3Mo4rDIf6r5Igs3kK1+N
BFWoiEhI/RLMpaR8q6O+cEg+XZyledso+GG8WkGFGOu8cLFZ+f2SHKNZ51Yc3QVDfzLmzz5V/fk8
/nnK9UJXD5q1B01QmBgPvjRZ7o5TZHEBkXJ8zMytkevlo/tpXkdc1aLYhTi2mZ0mI8dgwjKzmwHE
/FtPoURlsNkQsNvLKS3I/zV8pMYnMZhYRYozJrQ9TAitV2bx4a43s3ucU+z37eP9F7JwZQc+8M/+
453pM9m1rSMb80PTb1zvlCNlGFcqsplxBOOlXYVHAeOG7bm42h0RY6yRV8iSBwU7bwXWMg9T0HJM
kxL8fM5zd5BkyS0r8YUOrff/GQgNdRVFgA0zvMYtjR8DYhBITroTl1+fLODpSg5Rvx/EtprOiRMA
Edh0DDpKKjIdcpd0JnXqgoGuuErvquG0q4bBkOVTAQ4UshwCNvrJnwpGc7Zl/qfkeQ1jAJ5IPJr0
+fsFDDzCXCDFWPEv7M8jWGZwWBu24M6MRrIPYOsYbvuVmaWTbYhxs7TxreiWiI/KrhBUrdF/4A6R
DklBavuAMjyBAWV61i/bbFnVagCReeToL6WhoGDGYwQJ2tEcSZxGi3zTVtzR/AtBouLhc/Dwl13A
b35zJ3GFbtSeoT7p37++16LIWp4+klaE5FfxSz+LIbu/ZlI0ElxUYFJNeFoUMdCS4LtLXy/4SNfJ
d5hJrf2V6YYW+gSpxAgfTJvhJtACpoK1OUUSPYDggqK4y66wNi78TiCzmvZJ4WzLwx0JsnYiQ47O
uDijHjnfZczZoV0BEUScyNg7nFXG+52542GtEVuL8jFdQKbzTOex5jE38u/gF5latMWw+CS82DR+
ioMZ92m8z+jvjgVrlDx15eo9F7+jvTlnJhXGR75Pz9cuz25rRjUC1N9VNj11WWEyoeOsHWB3MZ5c
hQrd5M5Dt2c/KrK/UOgSBpWclBp6mF7oXZQuObHRs9XyVOjQmK4p52yB7v1GdCkBpfU/VO57XBJe
w1j+wVF/aWVSU0GKjp4XTNmqxmh7zmhe+YpeUNNiSoSy+a7LFUzDlTkSLeqWeo4h/ldzH4POwqUp
GQRqJPD4/5eBfbBCNefN80IrqlGahPz1f8Cs0l2m00gnZPNAzfoeOTeNsHGv8XUwvxEV1Ra2augg
j4cscof0+x0VXLbRPdjFF7RG13y3Y2fOK2viCQIizPA+3QcrlWUTHvCKffzPkR5aqNC+rSJTBgJM
39JjP43aTsRFlHnZVUKFNBrGT8HonpkYJIeGB/r+S1nnnXaTzjgQMBgGxPC/iKaETrB5RaRRd0tM
KK8x+tlSd1IU06qfDy7hKt3j4ORYdJr/F6cE79JBhewjiu7WpVHMrtC7SSYO6thGNBWe3iyI+xp5
iuKeJxnXDzkiPXaXMkZ3BxfcwMIQohYpoUg/mxaBtic+X/awxjpGRtwevxuWD0zfhHF91+8J4X1W
2/yO4Sti6AjEZko7Tt2Ofzbi5XKCTCLCFTEsjOVIvtObGdtq+fUk7C4LHFPHzUuply+lKxSJ7oPF
Yqxt0pxPjd04srYqYtXARIAITdTIE86DQ9QiJACC8ZymWnkwS8nF48/TCs/12phpVofulqAePaDL
TgGCk+Hf3rEX3xSGC2OFfDell1ksXdbfXn9H6oppASVfVXcZP8zm1xIZsptflmUzFe9D0EkTCzX+
XNOQE6WfR96WdOfXKDzXWZ3C2dnvKZClDi6xSP1dCm1SHEANO/0iif2w9U5hkmn1mxFvNxTce8qi
LiXOEfM9Gz2Ys+OweuOMcCsFN6gbp+VvKe87kHWFFE/2SwNMkdalcxuH3oaci68TCiMHuJSlQ91i
9b/JLrxHrwFVQQcuLdP3E0+6rh6IfZIJplyfLDFQPD9n5oTacdRWNZMNx+Msnobk/ikZipQYhD5e
qzhF82bsROeprToWqzLwDhsoGK0xiHORfC9K3i+JkfVJVns1c7eI9b8/A83dbuSA4KxxiXA5Rv8I
cGJOuJ7YLJ4NyAE2k0HPWGU0QXojac/GOkVayums7VdJcM20qiLEtyBxUsiLzKwxmEJK8kLoH5jO
cFeAj8kpIs3ozggCQ67HQUTVl+5k8AkdBappCKTBtWp5AKIs+pjINztyc4dH+i8Fq72Yhl6wEWkL
TYTBBKKc/sZxUw879dVBgMr3fxMsc/Jf0Lb6qOdnOljDyK/7JFqi618H+wDKh12tMRTJqcl4/oUG
JdAkFEc+IsZ+3uC2KHSW4JSX/FvxM2zciPPBPCMlqujMmtua2NaeG9V4tm2q1Qpj5OvnsGywY/Uo
f5AQNlOJ1JJEOyy0JPTih0GFQNdrcDdFIe7aQNyRvpy45g17hhT+Rh8Qf5vSDC3jcG+JhxeNK2yi
WwrU6CSvhSPlXxtSsnu3rVmIS0WXFgPFYkuP+vqkPXnHb/uQfi2WnvSe5Iqk6HiHTXu/JLkDu7vK
u/6otdoXqJauTuOnTZ0XHxYreGBQaL0lpkGUOfP5xwqEC771oDgcqjZeTic6qI1qVHikfQ8mUVGe
ZcUtL4g6y0YUnx50/lE/xmNec97ioU416v/Wa3j5vrhg/i9cegmKb4XqCcV/Q4RKq4NbaEb+2Rj9
FZEWULafN81UPXj/tciIdU0THRGVm27zMD8OoyQ+7ouA89quNXcsTpJYBv7xD9qCRB+Sg2joSxtN
kNMHimI+SWTGqMrexKhaBqhRldBuXs//fr1FcPewt/yCKcrOGuy4fZZUipHO2lP845asuoa/vPBB
PMSV9GH0yxpqPh9JHmLp5ursBzmUDXxtIfHNN1EBOhNf8Od17AuycFkGyPh5Le0x3YvFkj68cghm
27q+h4ktvhXHIMnYEHh/6XnfVzerEjVPZvgX3jM9kU3x1eojurkLMVRH2hc/02h8VL79qDOghSya
8VCS4+t43fDU/z+wG5ryuwf7Qrl8jjMUzMMxJQ01Kaix+mnMaOezYrNGNqAddlcMZtlXpfqN16Fp
TrjRyccWoO/4/ytjKNLB8ltVdi0aujNMGpBXEXYA7+IKuWXGKkXZn1rdnyDCYB8MNc/gxVczO+EK
evcpapivmqujTuNt/SmoCbJNw4ky1Unr062OpraIFkDFE17N24cJJxatobscDP6xmGJ0MyjSfxKk
bL45vvD+wEQeAx+SkR9fsXKU5V0OOXuDBr6TPxcY3EOki/YUjTLYRk53LOpsP4moPPZbl4MDfHFr
+jevKIUoO911y+OXayg/iF/sQoURL2kaIgSyZiB1U1aqLiS5C9xnkDeP66wcGYGvFC2tV9YfWfSI
ub4+mkVQ+zaakjPDaRvJFf+RbHiER9zShEo4QB1niM5ZezHQHuhQA0YMdC+RbvnfSkQPy3vvpODM
UjRn5RE29T7essrmufa3DjF3a2ZQkC3pte54dBI5/j0TgC5D7JWepSQA/jpnQphPhQnXVfiMahVe
THB29Pq1YNgbit8H5ijvYW9a7jORmyCOqZmnj+0vAc6YDgQcf03KpThEwIXJdhUT7iyllBdURI5F
8VmL6Dm22hhDqxFQ+Iy3gJmxG5bM6u8tC4HE6BSrMm/iXKsX2+CyLL5rxYvCH876O1bcxgQfVnJc
c3Xo2RynR+Aweqy4Lq/4a4vNPY3dzk81L0lS3H95K4V6eueRPj0jHLrHGc9pUaNABKbqfXkA8M8b
E6iTWpj6TG4tGG81Yc6e1SlOG7NmbUkDaQ8LvVUclCh4Bmlf0U1Sq8lWM5IngaeFlS45vu5jGsnD
I1zSkTypXED3xScR+Cn+WO7RyQjG1AcVZZSkx8P0ALzmRGRC6TKoezQZXVWjPEF6+fb0YETj+/mL
sPwptUrQBEQAr54jJvTy1YL/pP8gMvxtuIoAyhgn4GDFit5gTcndBRijwElADiNetOuK0NdpdebU
80OSjDuaeJCLDKwAu7m/g/5UAI86Vmhvn+SLmWNAk4YlTiWVTiBtFWUzoTqm7L5mg7GXSVXzNQ/T
IWWe7Fq+7XUyFKkb2l/wE2XaiXwhW3AMW3REHPFKK2kLqNDoatiVXXfFOH9JMTIqM7P3Vg3hKR4K
p03mUuBcf9wPx3uPvQkitLwc+9b76yRlEEyzkR/szAyEd8eUAGvr/+1YblY6ly5wgamZdCnarEEM
C2tswjAIbjYcuX0VOUsnOd1EitCmxBbgYt0DVyLQd5N6u1uvS7tWDT72XeAwyJWqmIHLndOkbcek
GiXyXho/6Yqcm9TUVZmj/MiQUROey3d6DhTBuRjM891XIaVWJXZToSWTiTXinwgiXa9SVfnNEZn8
3IveewXSSEEG/82dUs0n1jQzMPuFv0wLtOA5JTqwyKV+RpaDXpUV2wrI9nh/9FkHTPiN5ZQ//a2w
kxYwIvoUSlgeoPh9KXnCLf7gLYB1+mcFX9kPuCkTod8YXFfcE9DtPF+kUDonq3thZA14QGcKSgyM
kZBJE0hK7qsxYGAriUcYa5c5Ed0JnoIHHUYmbJZC9l5Wq/oFhXKoKVy4LZ7aVTN/X0PpSfhpqFnr
Mnv1gVK7KhircNkjk1G2md9lHntd1DJqt/SZQHT21/e9Bj/ExZJjOdTiCGmYWkq+csDHJQ7U1l/7
O9yK6S90GWgLWFWNYT+PVFUyl+BJM93wQOCOOzd1onLRjEJ9nuv/pXyQQnPwZCDk8QY/A9AkIVdB
rK06Lfrc1UO25OrV4KUNLIEvmnK5ld0fk8XF6zGjqemd1mMMDY3CAHIQwHBsjY6b/HTOUJ2tUOHc
o1A/l6k6Y9JC3otBxi1wCBJakVh03Oqw758Jb9REPNaTHSngXgmkf8hslXlYe8NZLjCBNrBgQVy+
WCEv3PEKfxVFRydXuNqcCm1+sP+SELK0/rWVCu2sS75GQHrATvu+3tPsIMY+ZTJms0Nxlsn3QIkg
yb0E0mRs/C7g+PO3AQi1fHx/3tgK+OmxmIGb+UTuBAi7OS5TiHMGFiGfyIYose4xuJVZqCe0ua/u
ykt7Fzm0BHzLO2s+W/eeKwxcAOuJRm5iSxgcRiDYIBpUftX5AFAqwMiDwzLnlMrJGRDYxKg4QGjC
1svrB3JdQLiLCkxWGG7JMwh8t7wzjEfAyO7A0eAEzdkvOd1wPTwLfYD7V86G5fAzz9mEdI6ANXJI
5b/noqAohT203bbjiXJPzeqkzZbhchSDIoYsTgjzQPtdOFXhSWck7XdFBA3V6wJjKKaj7TxLJdI7
+iwXUSeOBKIQvw21ZGQYMFYNLV6mz3jPT+fwamRDqxTJz9Xg32LLxbKFqoZmxFtAvXv2nbe/rArt
LIPvU7w6jyBl7X7hd0FSFC3JxjK5btL9WkSIXLloexUME1+HpHpmbNNI3A3xCndMGo0aCeofKH+4
H3VZPA2p6rzEK8rqpNoBngWiYlXUbcmdGyy/JozIWll0gV5rOm1UEzY7OG0CJLVBLiEOGk34F5jl
HCwXmaIULfxeUmL2E/Dqf8qicK3wy36MKsXsqlZD9KnJYX8GumlW5mmFREHQKOPoHqvOun7o/ZQV
Rx41trUwAVY4kDLHfn+coV9Z22MCXoRIzrNaUT8sQuu95neMF4TPt4hfq9EV4sxDUh5qTjVkxZ7f
0XYsz/llEFvQUp0u5fyiPCzsLD4dpD6fbv1qM5Nd7Ik8tX4HKfVkaDX3I9Gr7CTmcdIO/M4Px3/z
LZO7KmPkgwEXF4Re2Y01LKwxz6hFG0PUNx85E45IB3NRjCzaBJ3wFeICPFxl+VKFGfZFlzfpcfyS
fhRUlGCSuYSBEXstnrSPtvbII+9OJKyPhheo7UGHWqRWXbl/F6OxF8FdyXkIO9d0W94QGhHHayO8
G6+Nr1vmaE99cDkAcnjrEZgI2P40uOp2OpOm/GDxz2wktRiNxxZqk/Q60eXNjdpBi3X09Dgv3SfN
1m4ZNmfiF16E0AmXWXJR2MYqtA1f5PbH0Hbfoi61XFBxGRNMlM/ZN2PJOZ5wIAJKsQos9wuYNk+e
mEAIxsTulx/kDwrviV7hhqc5DxF5cKXqlGy9Niax6rDelaGGxYqlc+312wpjC/5/YH/WrLoLYCFl
dORkga8OCyiqp0K/nF8z3nLLSmz7r9DencVBHJxkRbQuEuvdPZNlJDvKYECxUDRGbkiQFqTaQQWk
4qQgilV6dr4nKQrLWQFjezyT9o3T28VsH+eKlbcYeRPEjmW5EPB7XupgnagemTnsrNkB550GLH41
33J8WSNcsAY53cPiW/3rUqW1EyxXWnWdrjoM6/0U7xexQpe7b2RI08VZvGlJbGK3kREzurbwEcdY
tE/fnO0IJ6kIuwT43szycPYH3OpDWV1WaQmq5SwdpKF5wgNe+UvPIjqDX8nOl0ceWumisUuSS3rO
bhs2QUUlFrQqzU7D0RoKhrJecrVuCRTV6HBdsZUe7RUFgkJK5TJtJp/4o1k4FpWxPmo9wGHiPj0t
tPV4UFc01C7iRQ0mJogFFmm+fUYGjjp1FTLkmowoGZ4I63SyVWQOawAGM1TGJ0niwOwjRf08jWRB
uJ3L8HZYn1LLCYiaaWaGTNizR4jfIYdHKiYA51B1nghy/Ygl2PT1zXYB3qMqJ5g4GOSDH+1thnHn
/gjMlGAL2eIQMdAcEozPJ/N9rJpBWw2tGTLYj1WIZ+C3WE7UNseEW2eTQiWZH9mYCzEJ/QYymHX7
+Lq3bGrCyWPANFAMnJgGcnh5IWEkCFo8JampUKZul5VXRU+hV1jzamOOophSCHOb9y5Ou2ART0d4
MyBJ6I6qo6zRr42CGhWjBY+Q+FDCV9EtEJg35522ERgWVm1BbYqiLx6Yz/zEas4X7iLAuS0nowOl
UNqDkBGFeSmNYrG4Jo6bzsHjDDx5OyREIBHSQWfmfX2VTE7NKh+acXmyps0WSCSa3frOdxfjzHpZ
3fxa3O286zmi4px13S+i6BVY49szVRM8uWK2cxUVI4XPUJ7vT8eCHeZCIrv0PZWTUMN089d+UFT+
9vu/Jut3EXW1+pn6DGTPlCzRJZF0bf78jkUSPjWqoYweXu9rKsLVsqY1PFVmC6YwWfmYNFwA0unq
omic5iK9Ajj+kHXv8VdardLWKBLaZVT/o0cNofoVdj9zRhhVZS1ewUIkhhZuMHjL2jC8F5pIQE/d
gpP3rItHBUxuy6MAS52wXZ+SjzuN0b9C893Eogy/iI3IMnn6iTfA0pOZy9lkA3OdoZtNoRvFnqHP
TNiK7mpEttCMVwqICadZF08cgdMscu2a+7U8TSN+X5WXZHTFZfTkRBaAmqn5pNM9+cIqYDAinaHZ
FD7uSgiLYpj9kc8p024y+5BR2K0NOUXZrEdDEbk4hePc43qOQM/r7Z4bR4qomhyhtcy9ftaJUuJ1
4eFaz552nVIsioJQBIC01pycIeraajnRCiTeTc9wKFsYzayjXXOEm0m6tD2ueFtAe1cCsKnamFM3
9pmuoQChAD4OqyA/ChP4++tm93lq2DCX1XTBvhrJib3Mhez9LtK3h9qhK1tCScv7OoO6Z3nZhFbX
90M6T3cD5UlRV1Walm4f+kbdcsyQxivvLB4Q6/kvS7qVX8mqY+TzjYK427Ljubvs6d8f9ALqUk7F
zVul+MXXVlIAMpua+csVa7fq1oJXsiVxljPcsuJkbZssnN2yafGQdCFOalHdTkYqeIGrbLbeC5vv
o7P2S77m8l5/HxaUtMNfBOlGSTC7gRM7D2Jch6T3S7EEc/qZT67EbNVItIiXIUvgj29gfOQfWeiy
31U/gVUUEfKtqZd2Ne0LOOVl1kGLN/SfCiOVrBolny93gB3svTnngLeK83U2YC1gZQ5VHS02kx9s
qm+JIDMrGuhOY19PRjPmD9YcDs4MUEvRC6T0aV317YXGG9YKCCco12cJMFLz9UI+DemkZAmN+bH0
jPXKRyhJueqE5699IeNerEde6ndcznJx7WtaEfV6MVdViY1NYqCxe5n2jp/61lqGUT50r4EX3wnt
CFQQsTq9/ouWFiEyXRnyx7Y46Yvphh2mF7VJMVIq6nHx01XSzEl2wAXaap12pbf3+jT/xgCWnoX+
7tHJ120lKm/6OqnfHSa7KxLH3vdVF0FFtfMZavyd9HuHCPzrZ011UaarzfZaSLKGNPylS4979TvS
svYlQqEiO2BxzDbYgefeoOomVTPIKzqmy4+Uye42myWGY01NF9Br3t/7XJ+zQP4YRlRTm7LxpVDD
PLA+go3ZEzMMd2cLpzXdsgUUXntsU8/KpMUqonO1NR/iaU9mQHifB4xsmdSxgJHnyNLF304r6aqW
e+h80O5ayhyePNhDRQXw/9oLAO6cSfdTYduyeCoQM41SxndjGqjokupgW2izlAyPjaI2cbbA3qKf
MqY/P4RlAqR/IuhI2ABpJNt/A2uWXkEL4MIAcwaQ379XF1Vis/GWLPoF8kqk5B94h/TqDt4TUBN/
o6w2KkezC9AYbL66BFs8RJ71y27iP3EYLJsJeKPeXEaLbRaSQoEXNomaSa6ACiBcmioSWInr378E
WuL080seK4HcxbDJuHkdwH7WWCHTEXBewCkM05kKWxeHOBCJ85LtMFqTpWLJQEQ1hSLn6J0qW7jp
ky3LfwiXbexSdL1OTmIk1INXa/5Q6Fe5sW9BwVhyC6VplYkO2NZ0iuhI2CSoDg90I0j342g2mn0v
WEkYbITb/mQzcUjtVKUzPbQmFO3tFyyn2qGgSQav6KjEPJ7TrgivwE2N5UafFSrzm5GkChwelzsV
d9OSB6NuMAavXm6GksTAdZtr4vckW96MAeftAEen+ir/5VnX9JoWiYFuvDK496FZ5j+kokGIOZZb
qFVOVfOyZhiJAk85KWJjVyjSkuwJJUpae1sw0XqlvdvoMawQCSyVx/0OSBiSkPm6Pa7uQ6O/Sq8S
f4UNPevAb5I8R5YXBwoIDbHH/IyNZIn3sGC1iurEYHG1FuqD5banBHWoXgsZT+qcAVR04SX9YiWO
M6jiwnXKpOuQPBllGWG8cMTpuJbJxjX0Wq7WP2ZWiFsmmnJrZT82M1NGVBHvCUhfMq9vR7qRtwiq
m2cLbvWU5Lx1/f/485bAvQRDxBxke1CE0a4RkXcnGNzE+zR4AGnfRnsjjT2oFsijkhzTbWlNfDiu
kWFDUjUvCASnxrPCa8RoHEdGL3QXj6xiNjMXCaDhzwI6t1832QT0c+uTYJ3Qv13uGsk1+L37Midp
wFBiZnE3xie/LkDL0mVfiy/Osyw3R3li9eZJvh+1gskKgvtygOBqrYYWBy640Pxz684s22G76xv/
8dUCZLQbqYvu+iVoLKGDtPNm+L4x2drkqEzJUVdBkx7g4to1SbMfpzVJdAWY5srvoocXVFeOn23N
NKhWme4zPBYUNkI1ty/nnBskkC6+ZiJUtCjZL53dsAEAeluEAMYmRNdFCeMqyMuu09R6mdTdtHF/
Kp9P1LzAFRp15PUyQD97tUFmEwFzecJg32fH1t466amMzuuQQe4n7A4DrtQnkQUmjcpkbPQCj8hE
m76s7f/N9cqTsmSd8EJ1SDcWUiq9+TsW1273v0L6L78+YwqNRB6uTSW0nheeg8/BQcReJ2xKeQC5
YcxiblHXi3IaTATcRjq6b5Wot24p1bhG3qXpScYqd/W9wbnaD7DP/Ti0lKQ8x+wmi7cCSXC6a2cM
4qNXruSw0h8kLBwEJGJBxN1S1R0exj3THbV5bngOTDpNKqrLlC2m13pmKgYY6V+3KamZZ1RCeZ0u
kmQzLrX69U7IqO4ekK5E3m5lZ4hIFmNbt+AALq9pjDf3s6i5cfFNnkgdXC70OtDxMvo83D5/WPlW
9fTpt2vOW7j34Qt4YXzDgYrAopycpThQJNdHbW80DS4kdUIUNy2nivRTHoplU3i6ylQKTbbpJ8jt
NKTf21sCXfuaLSQz+hwDD0mAw+VwJFEENIJgRF0aNzEwvtyjNbzARHCKjZJ5+2Z+riLkYnRznE+s
JKe0hUJRGwWJQQhe37sCmjIgp3Ciu6KJ0uH4ZdTewPYUssPWyNi/m9vqlsvCW7eIOB4KMNOwmex/
Vgn/X2xFXvw7lBbCJ651N4jxR+9DC5dmw4SUyVwQs/0ulUqLezdGFLkmovrszjL33c5rTxMUrsRW
WmZCj3pV++ovNqo9Yv/PIFG4++KOqCS2fJGIo6rCS21h4HNnjU6e1nSN1xPMaxBB1GstXkcQdSZC
to7AyvXzn5vZVx/MM9NJQO2zAmE0wiBG6kEXsNWXBZuKpKHUhgzLSmh6jTt/gzcmJXtHczu8GH+s
XwdnbZ84hl8alOKJSaS8uHvGUr5La5BvHHVf5lbdPNp1YJpWc7jCij9+T7SSFkzMRCmb8ZWv3EMI
C9+TbEDBDBjuX3muHokSEtXQ/UzWCABso8pwgZIEaLfJ2m0ks7cjNL7ulDPaRcQolW9E+1qQAQca
YcvAuqoDhoAZ22SbXuPkH+7qfRRnNd3fqPYMCl7CGVehLHI6N1NTL9xPqXtjfPC1YqMh2MQjx4wT
RKKVv9rfoG2jjNU4Tkms6kDgFlohJ1/XLSgnxJkivm/IVfyCDCL7KKLV36ZnvFd5jbHtahe5IF4P
kLZ16tIoFJwIR33icwFHAF9d2vdmWu9lYXvTRm7g6P4Ru4v7+fBSKsOsTt9qXoldeIXAbiA4sKbl
CKcsNICADvWu9e9OIpUIMuD1fqouJ0DaGkI8/xLze3BXAglBBIw1USoj91Iy9QG6+4aRaGIPas1V
E1ZcIcAazKWnHTaKrjYXz3pzGaoFVA5R7voUvEUFzSHuY84JlFnjzNcIbJphkGkxycVjJSNA+YMk
G+GUDRxwFx0ji5HKA62K6NG/5Y9CT1Ck9S91tCYUSFOKgUsQG7iPC/KeIEfta3e6AiVVLBwZXHhX
a6COfudy8BCJLx92ksdykuXD85jXo5tMBvatN7mVePRJ4DCNOGI7j9sJ1BcrsuZhmxyPZf0rtbNx
/URrTSKNuhtso2hEUc9sw0RjYP9neE2kDcxpIvoLUNO1CusB7lkbBeHL/z6PV5JDov83lwQLXk+Z
o8QQIOTl9ARJwzfBSct29/tV31r0XmIpNF2rd+x9LlICyi2q6/f7BSltVz/V2e9SU7s1fczuLOay
UShfWnonX3BA2u1pbd5vNpgFdWGHwH8azUJp3uxKkF3QddYqVr+X28VkIMGsSfavXoGgv1C2fvRi
hD5UXcL9UnWJ94c74g435IfGGVzrgUkvKiN1v6LYYSdbpeKFW+g6MxCZtpu24YC9HS0zCDChVBH2
PRfAHTbKzEfsSUIYUp8plFrwIKZeYnIrRpExXS5pjIp3dcyznxfu9eY3veoOgRWvfGKjurfnukhb
EbPEqTEyD5ik25nD35cZVyGg1la98a04ysNCdjcy9lIhj/DFSFZUR8Xe7NYI9+dlmxYlkJiq6G8g
4z61NkXiA7KAgNWUPwxLBAbQsups4aaWmHtiJwY82v7fxru/hiOxlNNa+fe+uMtzS+BF26FEIKvp
5vmeFTw3vJMUUtz+Xok4r2QlA6lj88iMrIF8OdQXpKF4GYY5qBYYYko8ERkmkizPrm/caXL+Lo5C
2Ttd6LPc2kgP7L3yGF0sV1SEFCsHAQ7SL4/jHOa3Jnwv5JaGSUtg92aGf6kO1NCrwXKWFeyAdI0Z
Nuuv+rwq2iArldGupljrEO6s4JvbxY0cS1VpFFYtc+UBL5sQ319HsQltxAWSVWSL2EHA8CDkNwlr
THE1+wEDOdjfCUfBovFwV58iHo7np/J06m65ivevTXM9HND2OdvPHpbP4h7lf3esF1GLKniqNc4P
nIAXlqZKcq7VoaWthEWRvOxqHNVTjkO+D51pt5V0I/EtQLemEA8aMsK1hDcjr7LRhy17oAtlRCBv
+60wf7SCh2MlKioA7E8W9xYyRxUy3G+MHh3n4/7pq/cIp7V7swTxfHy0M5RuSbE4CIGRDQOmCG6M
cBWYv0AprohLQz79kE9aZIgMW53vU1WEX21xjrFkiyLRBqpU0uuJPlJfo0OOdkev4xqaCxxpxptr
N1raP6q0JShjNF+PVy/FhDLQg3LvnWT/NTK2Q1K2lyOgKqjvjjBMJH0Di7/ZOShfUEMxM+ZojWc+
avCKdEWrfa5x2AFSP/rx/UD6RLuwaNlY3Oy+A1qukp1rwJKlk9ywVAHaAt2309z28q7LQ3YV+yWS
6anSVYvdNjj1nA5/ayjYP6g6D+O6avHGJbRtFZOrRbcXAj9qXc1+n9lHVPs4oDdledMEnyyhlTnY
Qj1l9NjVAlGrnnsP2J01E5f09ynJ0u1K5rZMqnZoVqx4TQ1Q7oWaj10O/DGjpRU5K95NTr3lmn9t
9RZF6izveT3CRFBi5yQDNr+x7J6cQlzNmwndxoA57+EPREoxws5KehUpppNRQKijdXcepfer0aT8
J2W9KpBkWZjROlU3wd6z7/GkjzpOSNZAPS9YmJWNDvfVxcpBmqfCyw+VW8gVtstdas01jh8CHZsD
kswiCmrCU87bsou67AxjC2wrxjv59bLJjGbHdAGMo9YrIcO+bgwtlgAty4L22lCtp+BAOpjHrffs
scT2RPXxmSw9UrWVIYu3WqQXBkhDzX65398Wj+lolaEZeRmcpZEdzhWbVW37yHgqyeK5bogv9zzo
5irZjxK2zRWomPTMob42V4wx8fY8k6E8wz9tmmadzTXCv2tYt2BG4f6pCNtU0nluqogjMmfYEeis
0/T515QLpC9eMeJ3/Ag8g4XTFLXmjKPut3FcGXqkvkwgkqUT8vy9eF6hhKUqwW76aDkUddRdI/BB
dGfopiSKX9Wm6BTgdElnB7nzkwRmCCeWZ/bW/VVrrn9+qyeKs6MpWxubUYdBu0fV7NDfsNjcJZax
qA3WaY7PqCXGtr37ZmF6jUou8dIPg+UeJ9WCCjLzpDZzH/BYQVxUiFLZ35g6yQAFm6CpmpVx83pv
CuDZ1jPLKh3AOFTXyOVAZQO9tDTUIMZNbdo5zfEfQ4tiD8uigq9XIwvT8P0gcqdIq2+krPmPmrej
3axLuGFuxt2+J00Wv4Q86eXaGzFg0Bf/UOj0grYlTPGTSXgvYRqa7seODIYOjAkMduNQcDTKcBzY
GDr6mYmqWifbYEgKS2PfTk+MVr/fpV5WsB0N+BZ+YAY75LoYbePsTTiomd++pQQxZRXKWDrSeONp
NQATDsGkWvUVJQqhwMShdGpI3fEJH7mOy4+1txynAA6KAtlwYgwlkgTri/Kq0Nc/PCUE0WkBi9qt
BA67WOxm0hSOPlMmlBoe8kJ8GsKmO66gi5WKUaDCSGI1DzXlikt1zZ72qNAkRXGDPhQL31AwCI0c
xGFeGHfZrVXvqiJC1KTNxyPijcQ6rB9NrrZHzVNS3TnATVikia0QMyRID4Jg/6ArSwOaPYPJl9+h
l31qBQwQyBHeTVHPLXPeI2ZSoTIfMBUmSiJlzOpv6lo06x6KxzCJLX9WHNLLX5SJCga8iEBucDvH
ITBH0L8UrpEeEMmTr5kyNrnlItLsxweCHIdwlNQmweRet+FPMPgtvKh5jfI45qi29leIiinqe2u8
nYq+PAgQh3Hg4DEbd7zH47a7yPJ1nyQISJM0ODAw8bshKTF5ud4oeN90dFaGXJsGMeaeUqyuKinJ
qTG3Spoiw+P09T9cwEJmd3ntxiTO8hRq5vIp7nW/YDzQAwzMrA5AEm/HfJ/wkBgLmvDnpMIrETHW
FKjP/PJ4FJi8YQHkZxKcDTtz4Zb1Bm+rN9nve6mRY/HNk/5plwKSSS4HXpPL3KodsgnbLx819vFU
qkhhSSTBP2RG8ufw1KJ0EYd4b8aFmBox+yUMf6YNyMOyMxdkRge3EJR7V9wyw4esBZ4ccSEvc3S4
T/vGiwuaUlPJyESlNE6ealVKeGpA0iz6OPPessIyJs/palPRomOFAEvSzCcn+81u7AP2FIH9tsax
dqrltYThaqZKkwL47Yn1OSXTQZgY/3/ZA4FfOOXDrWAiDcDhYoA92Kv+pKUgb/zs9aVwOR3Al5Ok
Lq5GEbIHKRVVUIhnSrmWBZPPaLmucqtNncXYQMUFK9VInpc18bydZwQUFzgqYgfubLQpf2s6J5OT
0R7Nr4vhmTRbKtEbok3ayHcHZ8r0mSl+hwWMQHENhsbaDFuc0Vqysy9Nk7l+Rgn7ygP8MDCBzuZw
+PEGyPDOGcJcGnEgWHZMc+wEkt7sNNLlIPBB442KC2c6WMgtzV5fEVqDmcsIMulrw3ioeqNnjF1/
oBboUyhlL3uqCLveb5Whv3CjXAgyIOdlQPZocSiL/mgN6+GVInybrZVVjxie3HY1oqZ9sQ4+zW1S
smrlkQ+isw9IfF+gh9CnEfBma33uFZ1R6RDyZ2qMI8vORswULivH4dLqT2WEuhD/pnAq9pic1R4Q
6JzF7QSeWdNyF798YMLK2nCUnSsfkT/yZMeFnDvXRRd3Fhk0dntKuUPRmCYPQXj+idDlyB7T5n2q
1u8ZQBUR1cgmIrDfLIEdhUQyytGzhGqDGXZjkGSiqP8ZzM8e/WOMWswZcf8IxrswspVtlgHaHFwm
rDJuYUMik1b62wHSA/9yRTM/dgrLk30gq+M28wtUnZMeZ9Cbl+9QE0XOXTFYeGYJfSrStoE9RQHX
gvJCF3PHchJxffJ2ynfSQ4NnkWo+6DmldsNI2bCyVI5y0PfIIOaKUJxdjh3IPWEXx+qIaJ9ZSatN
CQ+CB6opFy5ZWT317qAI0po2fSia9Inyyp9MuoR+tGeolrCKBlTqKYkO1R1+0IzTbEpGru0JR3qE
5BtzW+ZWbwGT6WYOq+RPhuyP/3nmqlTVxHGSBRQOAl3BgjENvq0SRxLyM3uB/o5Iacrnm3/lj8Wk
U3fecfNJETWeEfgrGftokWuPO4X6vaxgPIbc4ek9sGk8loaXmd462wMaiXoau8F0A2iRENp+K2BR
aEsSDhdSaH9pp1wJYWvPXxTPTtc68yO5owW13VqMQZ44Iok+aH76jFmy++q7LHN4rJH8rb6xufei
c9WhRAtR23wgMXExbjmOXzdKqlrMVQGFtIM46xNmakWmipg1j2UhvI8bR/Ahk6YiHbLyOcfHYSta
xUGViz4CdKvVSmuNb9nTDvEcwIeJsYKG/2JLoO/bNHNk3gjXu9k2sp12KibTTMnleAk4nEvFk/I+
lZB7TFHGLW8OvAyuTc+LY75QRCpxd4ckx2XD5lN2RR1HDoD8X/icTt2W3tcK8hwHjvaMixQuxxh3
hK85TGl+fgp2pzbDvhJzB3ZGK7EZX7mapnZpl5ndJMUizP3AjgO1DAfL80H5Y6i4zhiDwN2y//PW
KjPJL6yssazYXhgeYXd764jsB5vZbtTDFHEhztnxRhGVVy9VTWxEhBYki52NuYlj9vEFwImYd+tt
VqejpF5FpzxV02tj8I0dqOlKoELHvbYTxwe+q8AEVyacz6Fwzd5hJUG+Og08NM9uESUjGABA66fD
JLS2dZrYqZ3fFGGZlN+bM317i4OLxglAi2lqxdZGvk+ToyQG+aDweZ9vUAkigxDNXkn7Z7tiQx9+
YZBTUDo33WMXsQbbPfmCE9puu6yJWbST5VZwYGrLCJpt1Fw+qMEdQnAP74JFEaLBavVI9V9DYG12
wvC04l4EkM9s1/Sci4lh5ZsyBsxcwFANwnmGB2DCyVJ1SrVExoVZ363h4cde1/9xNDlGavhvJ0IH
23GbCNpYoHdTr5kzAiwttEvoX0y3jHUOWCrJD60L/EQorDSzZ96LnhuS1GA1FRa2gHRrZvyY64uV
CbXDo2CavhEL35Xa94RsV9fnEItwv2DE/QJDcmYaA4C9vWe5Uk19sb0d2KMPBVpDJfD2DKF2GMdW
k1TU9A8g59aB5nrsLcoLxDzkiDFTxPdYIEqtLOquCagpVjIm8FHAqrlS12/pdX8d87oodpjJW2Iu
OpcEpO1vWplbmvbWame/6Wpp6yzLpS8IyYJuwsllo5km+2jYDv2UBCo5si+C4mA5O4fGVFElOWyp
9lb3jzJ2EEGbYQNCpnuyHzIQM+W4/iO/tndE1XHP97hYKwHXiIWb4n0mVBx0SQpwfdbv4c6Kxn0H
o21M/1oqdpDrcWvdrKpt4371J/VtkOh77YJVbY4rACYBLYrrLAvepo9P5bnmhSW0TDCs2A/th2CR
al7/uq7FPjT1O05aNUXBaTjFm05Hujg6cUnCDC9YHRi8BxU7jchxJ4Gh7pBZzh2usUtOhhEzyOlZ
nXS3Szk9WquuXJZluiDpCFj0iNAQR3sBXJfx9t0SwfT68yW1LrEs5WQIhFCFKjLAlZZbPSJohmSa
fNTsP5anG6XSzjli1lGPOI2Hya1nlRvWL/+IFN31hjRrjy7FuoAedj/oOxcCcUhvWVbVHwuMIr3P
0OqvvyxK7BADsQv+9coTteuApLn1WlbxPMhBj180XWvRUa5HGc5DgpjiVRYU/zpufLvytJRvqheF
iE/yeYBRDCpBRRFdg/ZkfWy7EqFtmEbuDITb2auilroBGatlmAPLx0CRXFXkxD9tSF9GYW8MKmXr
GxeJCjouJnj2Ej5jMGSxpwyVomYjKLeMVihWZ7Gmj5Praqjd40zwD+HU/3rB9Sukxmj7+F3Rx4nf
grQ7EpZaWh4xtCZIIv4X7oT/fkR2n3kRcpk3MDu8p7rGb5bTHYgc8CJvblZyd4PPW6EKLJsc80bb
3fUiLYLrLEvoBgoDWW6BZcyWDV3QTx/+/sbcylK03z8KYzyTUA5nNLHhNOYS5z8xVvQJ94S1qYXr
nJJn8LepxqWMpB54ZvvvB20tRXKEbIc5gL3aI6fL9Qx02L5FiPPhnDgRuOzW7BmAQUipJFXolIyp
5ArPPHJsC5uvU03NeQ2QnhsJSUqbCBBGCozdq4pAma518jFiRsgF1TSGps8W78RiBeMdDCVJPCDn
uF7ahtD+/z9Siyc9lDk4RSWgZGmoxfbDpRS7TqqJVoO9CA87vMfdbjXb+FOQgUoF3h/tzMXWLPdS
3VeVPPOM7/5kk3QF6LF/hkk0b4mQZnXS4BOxU0W5uLX2nvqATHzUhoqUtDlHUOSY9oxdDhzJXfAo
Q/LK+MlboGD7fr1yIDknE2m6PHzZ742JuyqwEy6WSNdVXTGTn5nrMpNWOExreVT5LzOqzPw1UDXP
f1a7c0aP2AyghK3MmGNVUH1Wyt2GdqfjLuRE5zY1ptBMO30ZYNAkT2vrS87Y9NhmqizMzakZ55RQ
otGA1yDGQDBF5LVGkqc5t+j6iD+Hd5Ybujg4qJ6oLUark4Fj5bvdvTiLMV92nwkcMB/U0aC9xzdQ
mLKFQGr6Yuhnx+xp3kzGOwNMhRbC3o3qGMDvOVS9GVz23vVHr+61PIGiT9g0FIs/1/MOJMGScNA3
3SI4hcfpR+ipiG8x/1xEtWMxRDLhz+bZgkO6D2LmOEHsA58UsVLunDM9JsroU8UacAEGK1toad40
VAGHN9nR4YJX2ceW66Qz5BnysnJ8Q2/KG2upw7QUYkth7Cyx/6fbGPFEG6LE5v0D6FORXc5Mi8YO
NDftvvNLZJo2uy3E9DBloazS2rE05HWn3fAbiOwPHDFEeCpFR2tggdIdp1XlpV8TeWsTvY2A67qs
wNSORrWrvqurSstNQtcXN53TGyHmaMgO0Wi1lqHHIQvigd9/HYIW2ogYSFcGjVJXEcCbEwyUAEF/
pGITeI8BDBcDBMJwnifQy+R+xaFz82B/pbCTf0pm5BNG32Towe3FSKgAyEUSP01ygvPSMbE2o2er
UY0JupE/cxNTTGKh/pDQIejqzDKLyXkYq+9yPkWrSm8x/AJ7fU/jwWshSzMpgdVA36OT4EDc4dHv
Bdpx9aiLxec3MGs75pMZEGZyiS4IVwXpjViKnnQgm+d5vi0GBP1GaZ0pzCTgGHCZfAUuXSE/FP08
gZSSQpJiXoQQhDuWuG1z2xvOOFDLFhQgut6pGe9D/MS/xpVrSvELQLE1SSUMpLyLVe0Kn7XwWLDa
konFmGlo7u/jVbPTrNSej38/b/I2T7lLaJb2H9ClK/4uK66mYWFywbJceRiZ2FSi6Y8pcfNt9gDi
AwlT1s2oOeD2BAhbOYH3Y1vcUfgRxkAsMiK0l4dX33K3X6ZQXyN7se7Qi11QLnbH3PVjgfZ4WVo1
7GiwPhV4WUHHxKcfiKXMUwiC0mNaXmVPBeWjUkhBS21WIPLwmxQty42FIATWAk6UQ4PtEovJOtq5
R8OHpj/fAXXJz2JDvVqumo5yasItHUxTY1Xy7XHwt3zWZzmUF70T/DaoycQVspRRyOWqw2nnW8fe
EwOYQGD88Ymf1jwvSdnIaKr+WmjSfGshaOujd/MxfCi904nu9fDlX0/0uOa5tPGm+9B4Fk0sZxeH
UDHROIOHUOB+q2mV72+znRZcMWJ9heOdOdtQkwZPjLOY9qvR47NU6YnIB+o0lO6DGcIxasUGHHGZ
MO1TnfykVAJr7wZFWoQVrWXnf12FfY766XIynUEt1lfZKT3ueOqUQVogK9P0iIgitzEAZsykR8+H
X3l1nNtTXgL0uR1N9rOA7qAbPD0mmpr76YWjU/1ayQL3ORLdDj5LLNx4iWZ51rB2UNE6IaIAN5oY
RaXVPe30xxRBjv7sqBNUt8fmALIPcP4I1Nl4Wx1X9fsZ8dI1S1+EFggVgyhlJXrKuR5CNAHO8BaL
YmabAj3+/mV2112E4Qh2POLn/nHEZmJ0Kyibx+qik2vULIUJ9iYn86fVm7OTQbZdPdJhj6dQi3MB
Ecw0QhBk/VB/9/gpu/TDjjwFbPOQUgqOacD5Fra4kgjGgcvfwQWQVQvupp8SDnSk162tjPhJBL+H
4ArAUGJ2m1XG2jVwPHRnYQs4mUg1qCx2cMNI2Wxb2PK5lYbvPLPE4XovpYYWkRiiW/2DMhLm2CCz
D3iCebzI6zbz6mcBsiunsmCQLD1PsCjVyJP3ZqXbANqLV0OMGu4HBVYAALT+GtEO6Sq0vb19Alr6
7eB50PXvUxu7utJGo2hkFFrh/sy7W3R4Q8likuAPnn0Wsvq5Y7vdLcZXkoRs+Wx1EUvdrqx5VSKJ
DBOmyJu208yEu1V9bfglLwIcsjAv4l+Of7WIXggdjyTU6MfT87Lq7Qs0nAXJ/+X1Fv264nNBrM8V
C1BT3eD04Ps0MvUrLIO7p5WJcTEPDrEsxeytEHNR6j6fzf4CqBiT0BLhoiAnZJQw/10Hij5Bmzkl
d+UkMgdHKZKJ5xK49VparikIq4EWbgKzp238V/k26sE5QxbgQwLKYp1toVsfpHXVn9Q6LCIqP/M+
an8t/qWtiGzW6F6jJn4q6PLEzqlk5e+rhNgJZNDUCCu70KEEWSR5UZeMpq+kimraHASwZGavj2Qz
XUVo0dwju5wT1N5ovLC60lsjBW7AIYX+oc240AKPg8e1LSkmQmwYubcYy4iyttmmDafYu2S/VxGF
HWNbgxKJaY5/SHM9b5+a3QuDGhDHrfQwBnbcv4/gUqZtPwCbhalPZKzjUdCgKo4/F3Zn3wWwdVSw
7T7Axueb5qga3/8X/dqL6UWEb9qSXYxsloi9rPqcg64qRUKxJJfcdVccV8ViYOJfy5Dwrn/iPiYQ
X9IQcAaZ9rZP2bNIh1tDF9qmOkr2SRxBVhXIjAIlFnIh37jbUr6xCfMXiDnfZe/TXIN7LuCSCh9g
HA7wLTV3pZL3aRTqv+ia4s19KYMmAhRttd2H3CIrAKMuT/KSdb/HEMEYF5wXOZYN+N48kQLk+yOX
D75YScltZrhNPe7Aa1Mpo57jDO/28xWohKyHRZ9jwXw48LxXyNyORS/qBXS5AV+39ebqndepmb17
bW2W+w6QYPoEBnc6T9TSR2Rkmu+GIVxgR+89L3Nn/I+9sOGT+MmOC8/sQURbbk0RIs753Z/0WlkG
cAqPDVs798zFSoPXB4qqa3ZbfC3AWVN54TAvar4eKV3rZGdxXfEc8YM9K+14HjN/xiK53Xg3NjZf
6t2O/33rIBhOlnGlJG8hMwStAFH4DWzhYhm8fkBcqgEdSEMCUK+NEoodvUJtePat2Zf+gy90ajbd
fpNzib3xfiGonZs3dgBgJ84E0XskmPZFLMq5xoEnPi1bHKoyqEH53D4vDSlQORlGfQiuObOvtZDH
p8Mdcl4/FeOcWh+J5Fxoz6vGz/TChWbyfLUJqSXKGskdAG7DUAoYy/V1HPFq1MKvK77uLEUZ1zJD
ZfPv3Ez4ECHWh9aLcX35c2nkuSCV+U5CvMq547A/0/DmvkKtDHzQzK7uZW4YzsQiOcjPmHndFfry
Zis/kj7xWESx4+wREu6JItHu4WrDFVS7ijTLKfXMPrJZ381oOg8xa4MUrNWGC0C3BXWUtC3EaEdy
h1S14A3ImT4slv2Wf+0tTexY1DpXmpfcbKYw11Cr77ys4CsYDuLy7zUlVTchVyOirymPDAkiTs5h
7c3W6odm8akSKwUpib76nxSyv2tIp5xmA9BY+7kqJv7bFTfD20hzGM/edBFcg4ka8YePq8VBHJtg
ACtj3MMAiVOslCgDurRDmd8Zx4XEPKzNEbmXON5HcfejKmkkc9eMqXXQGSO9aEkRC/mm9MKkhx/L
ndUc7DHRAYSkq+zaWVBmGq7w/Qu0EAHYMOs/u+ZJ1HlUvg24I+SJy1EiFHxIllW4VFdTuuY2qLlc
1xBLBAfZVb+DK+jUsbJmn+Aedc66lZINoRIdlJnM67PpcCgf3bf2A7HdMIfYL/1UEh8nHK6MR9m9
oU6opFAY6sC3S3XDvMBoUMaiAjdwLSnkSj0+Ehl9tc+BYSQoUWtBNtxvIwka/SQgc/LD6RFxZ3+Q
gqp8wLOkp+/kLbc19W9POtgIm3EoUhCx2euMCT0DvL7oX8fDaiOm3xHPEQgZo7R2t3eMGkXmBUOn
2Gp94sagCCMjSzy10eOV6YiGZ9BfDUDZ9H2GPuKsdEBrF6bKmAv9R6YGOinZwC+dPbu6rFHRRKXF
0sEqWpkXVCU1GgAlKDXrzwOctFVNJuk5xmhM2dYCraeJDWHxdcvj8afuWq+c2frIoddhbRcb/qkp
MFyPDBV0BK9d4PbDi6Y4P8rByVUW87slAnp4O+X85D7diMPKRQF95rW8IGNRkRf8aMfN9Ac9kMoe
2Y4Yo8U61JQKNeNbuYJbYqvQNXV+TG2DWT0yXs48FseBfTorTdIHt7TpF2Vcumhf+mJ6YtUJCKt2
Nj/DGkxMQ3EtBtSgCgwVP7gOii0AhXhCoObwvQj6Cxk9G92hK09+g+qdK79mqWBemduAVlseROC1
cYQ+RRJVdWjwVyYyOrrI8bYU5XdYvN4DOsbnhlOfMMu4nAn9MOLUl+DC6v1RcrbClIznjibrDmD/
DeXEMeyzbPp0g8T/EEY4c1zSgVjRi6gq2F2qXpdJQ9GPbF8K6pB5gYKnk7FPWIxPGUynK0pGc8yY
AALNQQyKAlmudN6gmC1OkEA1/a+tr6BN37NTrhrfuXUv/+8wiDm7XzyPBfFoejlTXUNt4XhdihVT
NJp68+WrJdKH1xsrDt9M8phs6HWLr6Ja6u0aay7kGkEbZXNdDVKsi4S5qMM3pNJmpdmSs/bFUOks
7BQ+AjOAqXQATo3TRG2PusWAs/CdDm8CcPHdX0UapqjxYhLKtLocHSzBPXufrnhpFwgbgc+SSU4f
Lxh2DBRmFpBdPpx3RG72vDtZIZDwJ5mQPhGvde/a0z/+FZdUsYvBauda5JnXv1OJkmRBUkgfSQAB
qKoNZu5TpxHp9FJldaChtmuP5uEy63o+Y4wmS3cjgEq+ErcH5S5bngWsf2XDzajC4Kn0qXgFDQ3N
WN6u79uwl5RNs6W1jlQBg2N3jcdNJTAaVW9pwd0o9D/yT92C5gjyWTHBtbzZHRUWZW8B7Mf7JrsP
WMTZKfJiUi3+pQdkJ0QrUA93U/7uwlacKC7voAI1POHWQ9z5jYrA2ekO/zEXJwbm3I8q5mZ0FGEV
XDSX3g/TWAAy31L8vo+lj0dUlOqAp7LNYzjiHbc/xqQUJ5oh2jD7EATJu3kfLZUdlC0A7L0JsYWt
z6GJhtycPdump31myYwJK3TIqA3jDcNUML3FUvF+ucHQ4cyd/XLLnYRmsfK9lokDhfR3wK2AE6pn
TTAOMPNLeT/abkxTwXwPfucGWzdrNGv+IvGklN3ZxshH/LZZNDPLVEy0unshuDYf5VPjR+FdVoZC
0zKvZy1LEgzpxDRL7d/OFzL243mNSWLm+Lkx+Er/Q1xDqx41goqhFYqbgOpacDnPzctWJEyO6BEW
oN86zRvEb9Yx8acy8PHOYlsGH61mZBoBPZQhv/W7+x7dEJA9C6akpWVlxyu7bdhFAHxbTZOV/Dsm
64zdeGHjDsd1Bg7Zpz3cK6U4cIsbPjD/0Q4Xuvz+cNxggdoqCxrHaEi5kVZP9G2oBv4LdUPKD2oj
FnELhK4q+uVT1Zi8VhBm51qbU5k06Et1p8Cig0C7efu1irztiHqOjhMdOyLrUITTjHb56o0RUZWd
YAnLta0mcQa6+/x+JWKwfT4aMPj0K70374DjJwsjNljsmQRSREAIvrBF6da11qfXim8MOlR4Nmpl
NUKztl7uX/AN0iuWNmyLPK0fHHkqxtAfANlLpzbHZ3aQam95zMTCzv2k5d4MYmEb62MQwocOKzvf
TZKgWmicTOhAbBE4cOKSeKECnkEuNgqcXwfYtSmfDgZ5xyQJvfb0YvYtRu3lSn08DKTvl/k7oCAp
+YlitC9Ytn7prN0pCAyyWVf6REFBZ1TXZo63NNtP4sgAkVtUxHAAbWx4rizAEgP84Uex/klBgaAD
ygZ7HDlfrP8BZO/wDZojDkJxcE0X1THEdFIucgqOJ79ezw8VGiKdJo+OzbPydYEDgYq3zlH/EW9/
r6wfa13YKMerYDiYz4fsBdC1x82n9oAsTnTZe7n/W1aTeR5kdFb3gMCTT0jC5IWv00LWH3GEZ/GC
JFPWe/p1isErlC0/LqTq0SphvowCglLnnNtdDSRt6Zmb9XaIWpAZyO7dmXk237a/gNfDE8Iv+F3P
SzN5YEA69/VkJ0bv/fCicnnSw0PuG7PWtzOGYoMt/Rf3zdjBxvfsvza+KsaNU3xqjYt4Q1lxn68D
VQi7+OtCYTsPVaPCvY9BBe8XhWVBj2Gvw24OaYT0qNA01jtOg9Iu9dW4/msOP1zHqFb5unFoMsdt
zRJ4UcW7xVJf3LWnhoKHhf7T/z0mbpX/mUiLBGGqODeMJMcqeGHtrfY4i4SVZdKmh0+wSpHpBAHB
Sfl6TBzFUWY9/H5QB51cgzWLILKH5ibjqeCUchowXLJTFdTDzyx1TzvNVDfMgUmRFokq6mn4SKc+
IEZvFswBJqD9o2ft126lEt7MjH2CtjF6ZDqX71nzM9pkSnySbvgc1jc1IwIOHRv/CwTA8rI0zN11
oGSVypXKPIQ2kqySfXossMomMIqS11IkeRqaYxjZARzdXmDfbuaPBwYTcYZx4eYwWf02iE7+xD8y
IQgYcez4WeltfCskroJ4gbxTmm6V6XjjEu5OUhzwVj+u+f8tOtgJaXPRNEvROm6RSZbFNwjHPbrz
3YTIcNaWBJtis4eq8A7ge1zHtU/YOg4gNtAqEVlbAkdyL+sif33CA/5WI9OpC9vWahoizB4cK8jw
asNmD1i6etS8uvxbRdUJt9S8DLl+USXiBe4+7bRJUhn0bL9ECk2xWYGzOAjUHA7E0uUyXLhO23TG
2LaHf8+BnaRG3JjX5Jm60L1aOMJFIggrrH8vgGKC7GJUWSEXRydXHvKsG5DdkBNJ06fzYiw5cxjH
wClPbR1PSE4ajvG+KmCsraeo8+Shz1GjcXFwDlxHRBdEPx1YobmVtdpWmxLLbjPaLnA7QCfzHyKk
X+m+jzeRBLM/kjgyyyYrDrywgtKYMuG8x5lQYL6roCMVDvHRHHNizNBTNbZMI/Pi5Ggdzs9UEtdq
CVWSG5KgsgDM0SRBke/ep50gGtrgTvjAhB+CScrrP3aUjvbhyrBZRrdiEEcaCi73IXN2lab6SEez
ntHLlHQ5U8RVUQLEPaYrj2URVmrb1QO6Xl7NdfvZKSzTTZB+GAvnClE0HCceNVYPYimPhgmAkoLn
FU9xqnEjVJiXGNNgqzm2eLJYgdjToPGpJqRWAQ7H1RyZuoCKMc3djiG8FZ1PTM7Nav/6IdVwPXXl
GCeZtGtOue6q7zRnuTJIBKqrd/Y0/LNK4+PTKvdQ4dPm7rzBnwLNLSfsGYtvF9QhuKYSfX477DZJ
L4UTY7SAEbN911gLnBFeXqwOTnTo6rhYPzHotCXCyRzw16+qYYojaZyKxCjJC//ZOS3LEm8kdGtx
jyIIMLDC8Wan5xMbCOsgTG5TTSef+TrWLZByVktwWrgOQ3Sp1++SN6PraqPFtWXW4IISHIKWf2xy
mm6CW/xAgCu+o3p2fQLcgZfZDOscYsemt6+V96bdUT8Ip9nZux4rnv10MeOI+WYo9ObLkk8Z4euw
eRyewCzO0PTg4z2mJ9WiLpW/3HJBw9vjYDMdosq5ozQBjjzGFJt1X/s6NmB66kKlvX4Qk04KIiv5
KAT9hDAVtZT5FAuD8sE0n9NJuK6HBhFLcAg1b/xSywXNO/DI0g7VQR0kfotEH0zoM7EcnH0Eh1xc
0MxlchawN/8C3gaU2GXmH2JpTqzapbv5xEcnb7uzgxz35g4U+9XMg35ymY70JLZUeUDniwRmC2Fx
YluKk5XaLPg9LLQGXVXCowW5bL3jgRjSf2tD+B4b4pw0e7GkHnHwI+7xDHISbrgT/1jJ3XEiBMHg
fmy/nry3KnXtoPj5ErGOtGrTKHX6l8mNLXztTadLGX3JWNrl8biYeDmEnxUZ6UxJ1WPpjOoAImdk
CISKPP+BaaYzcI8qkwli8YmjUqkiG2Nh0lWoZDYUUsuNWKUoHUGubY260jYRQFrmPzTdukxmhukt
1g7FLHddfnbANf5Pr1gt5tt0s4BA/QUTRni+o3r6lnc4j9aDU7DBa0qEiFlosmZvF24Tuhhu5uUc
i/au0/PmkziVAlYk+jdIcXHeevFGVaDe4ODFMOvNW1Fp5TOEHKcY4x/OUbWVir7ZdlQmmzgtZm6o
sJI2IiyD7xlm1tkK8zCmoeXGy2pThtgloASksO6IeDjTQzrAZ/IOGZdbm5fmG6Sbl61PjMI94Qlj
cLsyga8z2LUUqwDJQu4QVMKvB75XVi59YZKHg8tD0T7UhWZelWuiqT/lEJ49bhB1ELVGfmxqFnCa
XvDZQ2uSy0x5po2MPFU3dh2pWeBPGVVVmAO9M+lDpXrbaCDn6YmjAVpxHDj4kQEaRSOjVxdzfOoO
DbKk36HLvqnvDR/jfC90dN5icnM440PL4fK9oOGETKwG3WP5SizU4WFmOSm2KQ0JCKYC0lc7LWWc
zPd73fliK4NlObBNRecqXDB62RmUb+G2gCBfjXOd6XnE8yS2HRYd9BwHdiXB42P6Z/ixcmud6lML
sZucjekKzMJRBP9FhMi4RY9VtSyMaSxOTweDGYblKP0aISYRxV5fd7nBS32mWj9IrHLvpunfFgo8
JJtbzuRdJrmdlZZ47/rn0oUq1Hbk6MVG+6qg6QRw/+mvAZc++pIRm+jHnFPGtjk9tN2gxhaSqFn1
6Lj2gK/nKKgZlUcYdQBOtD72GrNOLwGzVChCdMCWb0P2WATC11wsAKtwaGGlLav9F/DJtWwQRfGq
Jv1syBFOVi9HhopFh1dD0XrhxcJJushBkKJSTLdyfQPPGT6FU4WEYOsQll4VzrujUqwSQc4ZdEjN
zljXcWTHgFHNar+LZyEUicKpnxvYQSehWsfiioI/XIsmqJUIdjzegV8NWmYP5y8eG0Cd1zs9ZsXB
XOBuGaBNr6bVxkkrDAksrrlcAx+Ik3mLRbOAeMJ4ufzZk6TVSr+e8wlGrADtEfyE5n2M3Jqiwo+a
wt3MaLJdp9vsQfeHv0lpDogGNTQI0JGU+/wNu520IV8fNA8EjqNXbfsJjpjdSGxphZ39pMXts3AL
SMWC26dqINwGz8IhceDGSgxXubYkkUZSrv+DSlXfHZXH1eI/VcfV7+o2MdmpgWtxZ1zYXLC5zNR5
YxDg7BbhWFjSp/ONgcMRZZ0e6snbVZI3d7TS7xSA59njj4x2CzQxL4W05oCk93p+SCijuLtUgfRy
JhOCB2/6qfgBAMss1DNHNVo3BSkSuc55wlPx0YduzMmLEDTuQyDNCj8PhhFpJo6Bq5j9wrFlT7dy
+IVW9a89drFr9P3z/uI+/aqYkVsUc0mvRF/oJ9Sqmb+GE9uoDSIyBdMDT4HcJb4HtLn+X6j2H4R4
EmK+sB4QOmiHJkT4aTPSgBiaZlaUaBLhx+O0HUq42R61NynOb8upC2CMLHKY4Ly8WQSIGfH5HNnp
E/5mwBX0wVDFCdOZ647AZSyBFN4W5kz+j3/Yll2Mqj1XK5jde8aCzg7ectQauNoxhorOlc0RdUKc
62LrfspBlT3F2vffTVcUyH+JSet6HD9vClJa4Hiz1KaGCXSLJR8v6TVm0hXqYCDrDfslgoYFJkrv
V1J+ddv4Vs+AofiIac8E1AQs0at3PFLlvjwkAjKq6ms/1GUqzhO4vwEJxGjiBu9c6PekDfU0UfL+
5Z7DjvCO4uo6k7C2brcrZ0YoAtJYZgKegQt9wHVKDSyQ7ezvQ8sTxHkNbXiUIm3ylG+ZMffrr0Wy
YpkWmOhpPAfzAaqyXi0+lWFldD6Yobx+3Qr43Pdqwg/pw4A58YOFD1e4G4tpboByJojVz/CxdeUc
0W5U1+VpQyQ/J+Zva17h1imFi5iGhPkXf3GIjL94XE+rwQfp2AypI7MBiSNapMm1uGID0K4aZ5ll
8FiZwVN9iafWNMegznDGAqg9bELE+iN3PUXQn7pUyubXGPiqqW9Pu+NvED5r5jEsavVwGwfdV3Fx
rZIjIRoW1oUD5NfAs1tNUwsbT0Nsyd4w60VjU7g3sbY6zEn55jLM3Xz1BB23g65XCaf3AgmjTlpv
IxM+IMfmEQ4Fma/jqDArI6yMgzbI1IyoagKFXBB1tykM7c4u8H/YLUZndWi+CHR+hcm49swumKcQ
uIR+C53v+EL60IwtBLVDcbPT9faOiWTo4Z17UAUBPE8onbTmOXGfIHP40/dK/T/REt/jxpygIwlT
QgheFp+Wk3kdQCzSI7fRUjRHhwYKFXIbw9cckbOzCnvpgXaiqlkZvtH5pzrKhDxD0uQrY7LvQHBO
+nf+w6WjKNtdKxef5CEezcNuL3sa5x5Ce++7oiCs9wj0yxjYlvn8pTQub/VZb/6Peq27LdKyZ06E
TkG14jiMD13ms8ssFG8XZtzj5zK0gGpFne4m8T9c4hE/sVnoa99OegoDY5E4yUuENv1js2bAfOAj
DQs6ZO+uruUIXYUYskk/cbGHbTeYJotK3TOdGgFgXdkfsdI30+BB1cP2uAJ/aWmpFy2GIsoTpYOx
sTqjHmzKTJ27da8R2kO0DJkPiW3AN3vSlbISaGsoZ5KXl6NzSEcfFa90jkBAfNFFPecmXQGiSM8I
PWRdulJQqUNVfmEhRZI8Fh8MyTP0GAb8G6myliAirhvh6Hwq5G1P8wpQZOZBqKtoZhcFYgF0fxPe
GvWqC7BzrWbjeXkLZ07yUh1EPn4Qtauzt2LF+ct93RgSUqF29OwPud5jvu15VZfPid9/l6I7PwDR
zsSxjY9rfqwklENcfwsqqc7SUbOiPyZLOnuZcL5hH8wGeCnPRH47YzwTvbRGYteckA9zhzdN+7R7
RYUEsfpDwpQ2Rl8fm4vgxRUHm84uGBfCSGkpVLp4eyNvTh6wvp1dao/pbfsB5um8L0anVkOIi/VL
a2BJRvTewh1SmIfGifsWKzcTOSLPz8iVbLzM7mwNl9iiDtff9tl4b7VsjP/TaXCjk3kKo5/dfT1e
ZNhNk8cEtfy52K+s5wD2VXry6lmxcKUFI123mOsDh23AcvBK0tiKRPZxOKBQxlXC0q+s0IrcWaDf
8YwsGlHNHLFsZuaOdVNqnfRqosFIAGw45vtWM3g7STtHZSC/cSylhbVR9O5liRPzLHOck1UsaGJr
7sbfY8i6hyiXRc41Uol+7iHlDaRqUECq47NNIKUhNhG49xTzcUjKzgzJfFZY6Zffovk5BsfottR0
NO4mf/l3zQxqeYCW2r6TgsV3zrJ7zQ8D1tKBlTvz7zCXFssQJJyq/J/d5EBRNaJo64t3NsBuBJq8
/FBcF9L255a5FjSGm2qZHf5zZRbgjaBoUthrTAEseSuEWNjpv9iR1cTXJG+oZRmX9M4lkIUpjLUf
nUTE4vo/GTbRogWQ+U7BkIjeStzwuME4XwXjpsfMxRUCMHZgt/8iPNcWhWK1gRPOvV49c+KWHXdo
vO8sZFC0GxKlLgC8xTib9slr7ZLlwbnvJWIjkDIb/OQ6qp/DDymARx+uga4n8nQjuw0ga4H5ccQZ
6D7c1IWGxtaF1maQcTT0f1mHeKrtX7GXVnRysHglVqleK46B1TiHU8aXyFsEjU2lk9eKNQ9BzbL9
IDuqzfry3m0WFSSepiKzzPYfhQmhEPr23La1NvRor5icqV2Ok0xTeWsYmFFN0iCzOiWVP/aXcPmV
iNA67qBO87xq9RvYgHv4fLXMNG61LY2T/60l7kXePm+y0EYGLbpthpTmtrDYiqS2NAvSwuZrMVyM
9PaGjDSF8718N7o2c2Co8Ly2ht/rcYhcx+1m5KRm8lOS1Iix5yCMGjVD16TIOXF3c/QfXrZoHJ6O
m8TnG3QhJD5uGMg2MgAeWxlI/bL5H1VYnvXGkePvi9pYmTNfJm8y0UufzZcUfffNafwO6RVjUThF
ttb0yX3y6F981GvYWplqofC3/E1NaJscNsTbdk7jqO7jr6jsqbqp6BQgY36Kv8XQt+lRJ4AKLgzK
suYamXWf8EMi96T6LFxWyJLH8O5oWLtKqnpQGQ5fr2XXsTDs95yIEf0vDXKHd6d0W4mvXXPewolG
jtOhsIzZmrgFoifYIT1F1kyCwBvNElX9RSl6R+j0T1LksnuNe59tTIj2jjja9aR0h/1GB5Z+Np0k
H8TDLX4WTeFXxruo6N5fJgqfHkZSH0Jgbm/GQ/3jeK2YoC7fRXQ1I4A0VCMpGUA9Rs/W259bOfLx
8uBjziYP4IncgfJQyYCJXV/kPgutd9dJKTQbkHJvAyIbO2ENXiQ3knv37yGpe2Yj22nT5+ODpQRX
17poOpY/wgWCAUHhKozrY9Muetn5/aNamhYHJ9riqddiwxN1Ro90qPR/aN5z4oB0TDtlrl23JXJf
R/NjJjsEo00GqRz/hejg9ovo4q51uuMIKBKWKzJuLguxenA8pqHmfk4/U2o4OSd+IngTGBasF+E8
1kxyPN4fWhdLnKwZF6NVVtmgkKOR47SADt9aR5t00oNeiS4M7brDLcO9RyfmD3n7mfGd7aHocgmq
MH1FzgNA4qN0asZ+5yeCkvmoGmCzi38xsCM1oxiPlVdaPaH/BDnv7QqRlDUNli6RvztpLYnSXLA0
TB3o+UAq94OuQlyhYpBsef3r90kUKxnioiybsqDtDYcmiX3Z1aqzolWzQU0actli9RGWI3W3D3UV
aCClQNL7kdktCLcV16JOjHecT1XOqNDq4gVP2MzUeVNWZWHEiRU7WARAFYgMk0tvxBjbYQQiynBE
ByfL0KL/K6RQIdurrWKCiNkG7YPBH5NdIJGQrnfDUh4xhvn7QsaXT4/KSkdibC38E6p1e7J6M1wx
QYplbBta6Fb7cLbNezlGYteTWRP0Gi9zYrxVuaf689Bx34Ic0KhWfneCsAK1EgTZTTLP+ZmwkL3v
QCXBOT345bS3h1WRtIuVvkQIqsBTAeUrRui2NpVNMlw3Yyfxamr3ngkSlcv+iYxE5zp/g5EJer6C
CyG1GvNpHsItGl931wCoGvmUF3GJRqWXd6D4FQdOvk4DuI1V+y51BVvhhqRoCefZE//e3wYhzpmL
MutN5wr/0bbOCgosoftq3pn2r2RX0ud3jHV6jBHI1mXXAU/0cvqRRQpRiQIGzVRxDG7HG784eZlk
8bKU4I4Lz7JPC1ltK9qUuehxFef0l/BGSavJzmCdkmGFR8dwpMTlHUCiXtWUyz12eO3i58ddmItV
SKhnB+WjrGvnA4cAhLi0D27vJNeqPSkK3oCAyDXAmAJVd+po6cWtEmnq+N79Rp3yq2AWietd9ED+
Ll2nYJoGn+/TXg3cUR4csOAEiuNNiuaVWwiRUb+XS+7LWUIapX4ie5jDdgQE4JtLs39ctxQokt/I
QcApIhbaUSQFdHJzW0+u8ZyYiD7r3pA/bIg8/Wxy429iK6IIbM0NkaXGqLj0vcROJi9nG24mPETH
43OQ0t52X5dyB3/qgkzw5phib26FbovN40KXe3D5HZx54rMNGNwqKpreg8KzGwxRKR5hpdMs/ecs
prKKELazItAeCu26pSyPt5SZMqn9+wo+NyXFGSp2WjKhOd6P4mUiYEfEfWZ1LKU1wcI44Pzotprx
f2IHsH2G0+pDoccPNp0+RLtoP1NCC00C/qrKEXvYrH3U6tReli0LmvbKSwnIF+t5wQrB51y8irPG
fgyY2WmEOYMJ1AtRO5M4bpFqWmKCZIwX5LzZbGiAjER9JWVpoo6i3X/Jbg9C5EzMqtH4cVyqH5s7
npXr9RR0HqRsE7fe/WyJgvZK0Esx1BvBgZG+NPjy/35wt/6+mAymmOTW33HX8SBoQBkTDtGIG1tC
1QBqxjE3Oa0pC6ZNAnOJmt4ZnrmnTEMm9nehLB+aPBHOZzuyRAMSUcQvjU1MGV1wXKHKG0RS07uE
22iMOU06JOz3mnpwqAToO1z3MLoBquyVWeFeUnfGoMXekFFTDo5Op6Xmf/kQ1g0FEdSl7h/Txc72
aSPHDYlh53LoI/RfkA1LcbG5WpitVwNQqXHwkVcSpBmFZO//m67fS0hZtHANjGXheWisBW98TlKz
HyBAIKU49BLvy/c01feGbvhxI4BXS5+66FGbCZ2XfYR7mgMIGu8ex3aBraso+1+Fmmt4ZYde+d2L
eSx6QTmEcT3q8M1O/xrFziG6dGG/BDSnK5e8FPYjAAhMCjx58a19JLbV1PjKHwGP6KASQ8onDNBB
vE7LFXWUySYg74P9xQ51/hTJTOHrlJb1NxlKYXvazU/wDz1GE80zuyNva2mpN/qQAJqddApFAIak
8JKBAsd1wO5OCPMcLzhEf9slqjOgR105XJx9u9AenSPLO/2ZJ8vU6JbiIBiX57n97xh1TDGZcOgP
/MYTH7Xd1js02OgaXMigeFNLogfH1IIZGp/jVSPOlQFgt6d4kjHm0QJy5T2lgnTOz4Q66GFCIV9U
80r6aZ+AeBeuAOznkyutJpMXa4Wg+asYNkPNd2jbsMHtW7EzX2OW8KsDROA+qR/2gvYt6NGXwLT6
TCzoFzDl0ZUW0yssj9j7UTNdO9Cv9CEbAwJ68/lDiSkPK13OAdTIzqz+vazSIdVyXw+wJDlojMxb
by8/evvE5xSrHmWOdUEex1LZtnYxRVI3YmY92yxZbRryVvnuj89t2q3jjy3QcjdO9/4GC5DEvvgu
Qa2UIwiZFfDqkgraMpy6s9A+XbsiJwUOQaYPaX6ooM1ZqcYphI9lcOpDghiOZS584SNcmU+zBGII
8GtpyhhILGCtghO7IrUV7zgGKF/pOwVbmiV1qPDfv9KIUzSRC9tZppWYGCdvKtdyD0cNLbjLPLJQ
OK263awmmZHClBKW5Wcknfo62QDksStY0yk16TrwXzZZl55da8Y+WWP4uvYxF423Xb1aA+Swc2Uw
E3FhxmD1cj6u2KIySynrU20KiWUUxRm8Guf4U9Jf/pJcr+9vDvdTbVueXxfb79dXKE3pd0QIMFxG
wCeyNA0jOwhq88+UcgIeGFHF/CD74h5EzWYN3wYqndanDn3d+n6b7swLtn7hCdg//7sRRzZ07bta
UphbvzUiRinHrQ6ynzEMBtBaoSJJKFWyDjeJimUZKh4tP34J1iKQALqxhk5l2BpvuaWmvKwCQNuF
4eyLo3c0yUgc98IOh2AJDDx7GtntbgMoJ8xefJYIcgI9Id8QKyWL52/O6d7DZ4Z5AES1J7WT8Jev
vMgpl3eAgRR74xdtW1NHmbow3wGjid69VLUtmQkuR6LSbcFA3Ipb37YLfQpzi3qdOoCJiNnW6pXU
0+iwyraASl4jinxBBCsUv7BK5QWeTjmvwLuV+GDZPY0ugPZ5MWpPSKmiou7qrARHKk8Q+8tOTTDb
Lo9/x41mvmtjIRv3wTQQhmz8T+NxdNIC57GPvp6joxXr4CLifLyamt/HWbf+qrhuChMlxxZ9kmy8
VElYD4Mm4Bd598pBwiWSStPP2EuVMc9ntHxQtcaz9u1laeLQhwtRhMSVqvOrEDAcf4k9og0Lf58v
wwD2z24TYtsXJsV8gV73gK0l6ty5pLiWbkNt7vLX+0etGa84oymJ1YR7re2HNyHNkLJ2UsFZvsrM
awsLskXblLsWOvpL0olKU9syUG5rXVmWObzYaKrpsWj0pM4ocbTEfgOO5vYqQV2jb2/Fsub0QLhx
elU1QHOv25ENSL8pGmlRA7F3TpYFoTQDFpHBZaweYWucLZ/QHyDw8DN38ecpWntzE7gikoVy8X7a
hj0rwBz7qS8xaX37jkyWlSShxckTOXRXmtmOXmawnSpb4awNzd167Eh8BTFT65YfkgNbcNeziRum
Ok+EKUosIxPjJTo4JZiBUAr3VhdQ7VG3J3CSe5Z/RP3LtHcG1Mchq+X5Ozinc0pvKGvhjon7u7xj
uGoi5c07Kop/o7VcUe+X+blRsU3kT/Z2/agRPz0ZgDH26An+XyxXCP3QIfxbJcLNQNl/X03pvmoj
cN6a0ptKXbeOz412ttkdg/bSpUI0FV2M9P8DRhrYKh4TWT6M7KMlkmLUrKmgOA75eIfIU14lj7dR
ncyQEqUrXxUJHEoGWxZH4wOHCRBMsZ3tvCIm/pbJ9pECC4lRNpOHvuO4srVlVWkJPn253sCugI6O
uJAobUYcpvNvyA8AQr0z3T7ZkbTWZFmI5lCYNXRbYTwHrBXlneCYld9dvEnt3AU295Qp6kh2kL1e
h8s0APr52k/BAyEGT8GAyK1HNCEbR0QcS1R/WIhA6khoEwJ9ZBNIcLUxSTZkQ9RMfxJ0lEVYg/Fn
W5GzDEqM69TIPTM2Me+p++uIRxgebfJ8SJgmQC7+/iZb5UEXPdRxhb5IZsftIuUer4J4Rmqs+koK
yGd+LLhXzVcRDfdbkF5cBAPS+M1Vna/hGbL9cE3tqz+yRcEky6XuOtfPSBEjTiW8sW0TzRd9zczm
HcNfAHUKa+l1lDJ2I+MT/DuOJHnwQeMRSBOT4mxzO2SGEL030bi+Zg94UkLmevSeFLvunCZFkoRt
FYB1LUpxubjl7wRbVMkO+l6ehs6FaCmyODOdP6YrkugYp9zlHDykcJ3TIaHDMyZhYrt+j54RZ+7w
PmRTx4AK3Ln/qmwnQFb7aeb6G5XfFP5xh73ZlrrHRNgFTWhRRTBZsHjPQ0TYYGqLhnFAyZoXKxtf
PEDIz4/RFHg7UYbJgSVffd/sc9PDepEZX/bLl4kN/Yi+m+SqqRG5LFgRiV99T67YYkPPK8LyAhTr
MhWP3m8vGq+d8x3FvEnHRrqLZIVxL5HSaX0dAjztu54DnKPz9ftQKZkiDAbTapgwO56GDkptECc+
IOV6ifX5o4CNtfxbWlHK4bOFPwWCj7sV+RbmEnS9ef+IqasyRVT3PewYyEx0leOiynySMDNiP1eR
E7xfvzc9U/8uQe4I8Ibnt6msV906KKoHjvRQT4ibi8UR0i/4aqLvR8pojVNW0EyvR4ms78LJehI9
4FA7t5Mn+xZyKrEj+yH/1vLzNx8vh/7hc2sljekkKu3K34lVzM7CyDjyLVeQexBGXvIKeV9gIgA6
8RwgEy1kyNaTzsLtUvm6iCepz9snP+F+hQrWR97Aub7rqDCdxecEYq1E9NZCTolU/piaiT39UUbz
hiu4VOCl3yU5NfJVKYp6E59fBrvEVu5Scx4Rc+GQz2FUgG7yofd0gsFdI67d4fIg/CMnnBmIR4zj
iBAs1lsLi47+dmi7Q+hxB/AcFouXbw+G6im4ab9HP9ZBCJyZ7JNkEXSNwUNYBUVCQYK6pFpxU1AU
tsxxxRqm7d3//FA0o7jsqK34RsbntmNUGEplX+9+LWl/t607yv0Q9GQEqjWHczzqgGFbyjSVuTdI
he7WtE1QgloVE/kS1wdXMIl36wq1/DKrdgrSD+1t97JHTbl9fAOjjl6WJtE12UWpR/E23elfhCMh
ypHFH8tDianrdVEhK9MCPWXPRrCwm41n7/gsjgDOV0lFLTyRY6v6cK1n2kAU6/ivUGE7+hTBBQht
6ALAVvlwv/hfkf/2WWuNb692endr/Jaw0VsiMq0Cw0y6QFMMIWBLDgAHT5aDAMNoFISOk6H5u5ut
wib/RrYYNWItW4cN6qF8a6zsj9CI66CV4VvilaoHURENZAAbdTbFtmfqVGWLG3dEW2/2imvPbeTP
Ih9CXwU0iqeGzMVEACD0iqyAX4YThLoIz9d5f8MUulmLG10yqj0CY1ZhVccSSX3qknYfwfUXGe2G
VoIUvC3xHRF6q1srJOka+JDZ5kdnY7ZPuSA8KTS3P7qVMi3gLqtW8pY+mztiPp79Jh3BsozLdvRb
jkaUTgxi3xCYcQNlUA5A07aOn1FalGN/y1TIgVbzcdGz6OCP87K2hXb/F8QXDhZ3AijiuTXyudoF
li0CpP46v+R2wG020cJ28X0M0QzWb6JvV8to6RqvK8DLWLLQxffX2ipTihqSG4DOpmVb5cS1TKbK
gLF9mV71s9t6T5JpKM5EJndre42FB9PGkSm55RDxNnBK9AH2uCvpcoiZEPAr4DiIFh0Rq7u/5B7e
QF7XOmGi5F6sjsrV2PoR8i6uF2IDValLG/wjUl1tId+phlTO8pCe5UAOhvk4NFVLjsreH+W3p8OL
JN4qdC1Ne5RpDW99X8QESEyOrVwzIIn7CQLpzHPQo7eMzWt3w/yuT/wa7xtFdF/0VljTO30O4fUS
26ML1t9BOQ6D/kjw5VTCHd31gyfDFHJ3LPua0+dX8z/EJ4i0WxSXRIpvo6HFwPawr/5fu2XTyFQl
b+tY8jI4BJG+8Wy2FYMirVEvd5a3IAvpJfLvdmUC6v7gmC7/ZwSqlmJJTpQ4JUBsInMn90HUjYLf
nZrx5j/xJH0EqUnPY1MbgzYPzvpb+ghJhDdgWyGR56x5hytBep/QtV3f0lNpYhrARGWqQBgm12VT
0QEXQf13jfCm+JhAGPGr7CFcsMQGxDJPJHrT0OboELNxRNnDu7mwLMWlxpK7ktd2pyO/V4mdQWNl
osUsqheoholufVLDttBPGBo6+DQMVH8i6dc+uxf/asizG+EAqDGw9Hpb8yeSlmJcVqFe8R8lh3RR
Zpw+zuvM20EQtzNQ8s4hjRGYNgIiA1ejKmgtg45JQrNLDNL3T52XwzuvPJTdLCcm3mK6bKhVotyF
JFr7Q2iy/t7r4VdAqVcSKNEnNjFgty9cYdT5EsG55EqiBAFYfoCRxUK/ukTkDaz5oVtickTktWDr
xMMQrdSK67WC4gHx3wI51KhcUhBVY3Gc0fCnIpuq568ikBY6gIExpy44IwVS2MdhFvzxU570H1Tq
0Ew+ZEwo3EabIexCvHeoPmHcu/qFDnEShudT4AS3N/sUckrBv+lNgUhDbi7zKra2gf8bc/l9Lz17
pT1C60Hgj/ZaFbGj4w45GRjUFpfu0hsDF0ad3zEhh3/QcEuQ5mnnimcii97Z1jM3siY1SQZE/pLi
BhBRBBZKYhLzfPUqKzfmcCp/YZLbGIihiSNG9FFE8hEeQtwtZ/tv4DrMg0aPPM1DGgOOeLS+dCz1
pMIyb4x5wsrHeOgQ7MNtvNXpUrGqCKwIzOZNeaiAb3oSkBEqcHUw2xq0cvC5qQgUpani1OV3UXsQ
QVYpU2ncCt7h0A87ghcHUC/0T/Zfqh9E3IXvnUSoPTsfJXfQnWrpTmb0cGhNb/69RfHJVy3cDRqI
OHug/Td2GR26sgvI99KmY/GVXFhhAV8cW89oofuvwAaMwptyFTwf1fnORIZFEPzKclM8T7i+AG6A
FBxaSqJ/cTwbNMjmqAZBlwiOM77FIxqMh7PGlxGglYBzSRK2WovWdEm7+TYxcBaLMH+oLDCzL1lu
bWjQXTLt4oWceYNakEEIC5UnRTgIgSGoBmoLhN1aEhBtn4Be+ikLDgRZUs+fT/HRZO2JDq4pRb62
keQScbKBN0U8lKHTuBrjeUgsfYfUCKYje4IlZjF7TDuTvIkIuGETbxtd7aAX9XBcNxd7cCrdjAai
NYdo1sNFFo73d+x3e1ZvenYZGRPrHwXekXdlg72IROi++1wqJZUCNGBcIPrx9zu6TgbxMOippEmX
Vcybm16uboJWsTjQQpcI7U10covLAfpmlHMab4cuHkXJK5/FX21N636VvpbtJwDXJHhQ5DcSgqNH
7uT7mtZq6NMfTqB06IfTtJYcTKHpc7NXf7UU90PDJv1BKFTX/dBt1qSRb7ldaIzzjIObNMue+hRE
yro61mXUn8Cto12v7kk1SyTB1zPHPmL3fQSm4Vig9YQxXzY+PfwxRtU4rAeOOUCvVIWI3Zmsq7uV
pvFmmZ7JGUx5JQb4S3iF4RfRyC5HQvhwyDnxpYa5rIlLAc9+ZweY4mOD/JNlo6pe6WjIjzbs0ucU
WgePE0LovC+5klTgmez2/3ZWgjJh5tNlEscAndTicrGLRXEaSWF4tZ4tiQ0TjASFfQEcCuIWOYaw
oGB7DvlsX7m/Zj49VuzB11D9DUNsRByzIyOjyEZEwm6nOQ6qXILWMZ8m33ipbwrM8A4hY70IvrUv
fuZEg0Xq0kKrckc8UXwFS4Z8c5bahj/FIUwI0Qyyy5vTWj/EI3F4wvJ+yFmRipWa9FIJyUJ61NYP
qHchPwytAEF5GTXP4ds4rSFShXJYRw6SNKcga2T8Qv/BMYbugLeHASJh1X/5inCjePWlRPwuNHtK
fa4orFp0BJfwE6GP4JMqsNlFk/MsGdhsPbJQH0RAWTW6dT76c0bH530Cw9Lwwp73vGjm8CB32xMb
D7jEuW23yiBNBPNGtvEKJ6sNoCMeWOQRgncpsS/ZiuzIH7A4M8sGP8MMHjOdDQp38bn4C0CLM6t2
nNzpz+waCaFv38ZosWkerVBMSnkAbfXKF28sgm5aEEmijEUuhLp/CHoTOPlZzsjddY0LB9CVhmi1
+xFEo3cAfYbe0d/lqs0kgzhvZ1cIqh/Fy0+dv31Mm0dGvTEP2VlOFX5oM7OnybmzCFLgO0MIwhkh
iirapM1/ogRctv54zHQng26t6pAUJBx+9Rh3unmVjr6wm4khYnR6/xVHBkF6WPt7EJB1vR9qfb+Y
4i9WvHenUnNYfOhaLwtRrImGY7OoiQfPNBZbbkOn92e32Sh6P/AgOJfT1Pi45UqtGSUjTFdbZDsD
97UQM2tdSpJu2unbeeEw2+fEPYLkDYMjAp/ntZGsADeMHyKIF6w2jZq2WCz8rL2anLwVQrXNebKv
43+7iZ0Csrid0RKKqUl3YKIjIYzcKlJPN0GL4yw8i28kN4IRHfi43jy8Hw7aTSspHtzvx0xXlcx+
Yd2KmCFoj7ncadSc4KpHKi9HsHiSdDhsPOSj43PMKIhzKYRs/TeAQuBm7cL0GnYuCVxGSKXhQn6k
MXfWxQW1EXP4sbjUyBd2mO47LYDPtS3KphPzRQNuPpMrWuzhZDPDGo8fLWjA085LAY8fozP6Nr0F
UFTGMycQNzhZ+wS5BY8WUNYh8lxm8RDVurnlncl0zCk3DJ22GzCf3Gjc53YM+CinIZtIr8RBOl4v
oi8OoM3K0G0rpeYT1Enko6tkgrjQHhsi2uLgcjrVUTt26phVw+FJvtQuAtw4RfDDqxIx4iH7eq0c
mCQF6Gp19Uhc+8Nf1/ptwK6979dcN8GLjzber0FTUcZFve2OetZjU4MXv/vgUcDJTQAoOTedIIjl
PBnX4R1nSpctpXXVK2ZaaWf+pSuS8P9MVDFXDKSPS17b5m2VXBRO4escTEL/c/z+BX1Ig3hx6krW
j2hC4ntKXHYPn/b9GKLIVe0Y33tEO1yR0XgbQpjL871pYP7+5lUNG4OECKATCsQlgRz7KH+bA+Bu
8vXM+bS6OYYXtUCA8VrwQosVzLtk1II9CFiDT+ej0BOLJomekIpC+UyHWzQ/6bmXSdGD5rrnarVt
eotdPJaZPIC82kY3095KmhaSVkfX9TjsmQcyXSpH3AZ56XrSKHgOC5mT5uI0LmvXvLRr75I0helG
68IqvzIr9Mb9iwpSt7sBkvIiqx+hH24L+wfZpX8BvAKSgSAf1DPw4nStpyelEaPdgRrju7bEeN7o
kCwD1nZo5jkbB7SlChY7culZvBsR4bbM1qWTJs57GLfIOcRszOLputnC+fTtVAUWH+WoEEkTuBMS
lEj1LgUe3o3WAKaXZiSML3uANTQkL7UhMaxS4+Ro/2jUkws934VBJ+DCuKES2bF6oKRD5lpf86Lg
8BfTiqmiwlfsrMgUPRH6eQ8FSM80Krpigphfw0LP6PCxnYcahHX/CCMMZ3cm0pmvN5ATB3jMZHKu
6te3HwSwrL8eGIbfuGkqRlGkn7tJRJNqx1+OvDHry+z5pq4j7mTyEjiwkP8Cg8oz85+t7CVbXPVN
s+isJKuhjv30oXSNNQAdwv8ndks2eYvXgyUqb69uuPJhTC1U0sHj2wBUTBpWG/HFt4U975P3U2n7
4xkWYycxfIbVUd5/oiANpuqUA1fEopcnrjHkN2WvwXgfzZz2CXuGFbx8Upft6NRjdSbnvZaA8U+q
wh/hwzpYSo19AW/azNifrxJixDFiAYigAzuUE7t+RdKP3S9K3mx/frjlTXlK6Ylj7vC0BHr7qhgQ
IQFILftf8wreL6ZWSKbGljo/+5ir8wn+X+fBeSqw+Cme6z12B1u8totgh7Gm48QcHHwqHeKC2tqW
roEMOGBDMxeMSa9WLS6r9ToOrkNC8nNsV0If1Gl234alIdcLBHpW9010Oki3Xf7ZS3vdEEG67o1u
m4eUpuvBN4p3gkyYUTj3wmPwJiakKksmD7a30K+jl2EpRAYEhZxzZZWS7DiA5BStacgC8jicqHTI
h+o/9pZUbkAy7jhZG893fUUTFMEeYGhm4QVX5nAVo+gLXWwhsWXefuydRqll54VaropOTHvTqqtA
1w4Zu7w1RVZsLMO9GwUFdqZ4JWdwG8Px11G0B7uD4F4u3AYiJv1HU0s2aHRCRy1kEh1xWjt2fqAH
GOM8StQloUINcFfTkWocQqnckFdyfoA/uc3PvNQW5oKaDkk7Zhw2ab+y2yQRqhs41gdcz1bF+VLy
h/6LE3XrIsfylz5OLYQgLbBYu1wMrZOVAKIVU5+MwtXhw8MCzSYCy30UNsQb5VXKxpgyoi05VDiA
+jrkeXkoFNC0P7wbjzA0XUZmXs92AG42766L8QmdjWaiQL8dp7jEgpGFypX1AQSji7Osnc2dQx5N
OpNYl4XScVSqTfoOcBXHDYpzPkF0AQ+/N2rHdcUdPxyrtVRw11wchOKfhTAPK1PLrh983KG9oV4K
ztknLPZepVG/Xy81LIhY3fQP6gD7rntxI3g1PfR1VnCQ6bfWiWVhQ/ADi9gD6v2YpkSagMBC8f7D
IOMHoXWnMNWMyWvwz5tYoCv2wParXxMydp13pEQXwmEgG7sbANrfXB7V3YmY5xp8uZJ/GwIC1d8L
q4jKNFzjPda6XkKJ0Aqj5GUrNSG3QbxqIgTpwMFVgbg7kYFDvKykv3kOdeY7tMGSuPyO/Av2n07y
sLg0ju2Vjn/PB2sV+E3+OHG16escAtQLS7mNtBYyctX0SMh6WuDcMJzYlLGE4udIFxCjjrIULqYw
ep84nCCOROmKQ424Bceqq2zN9nk/aJAyXEfC9GNmQDA9F7SBsE0ZafhT3fA2JOwbAuWmiP+eHYd5
AYW0cC1bGjf6Lsojz4OcjGoBMmDQVbpxzn9vfCqegEA0SEj4sduiMFKvaSi2Ob8UMsOWttncKkGu
vNDjYlwFjfJw4ntYLMlO2kQiA+qjY+/SNuaNKw0uK0HhO17Z3ouY0XFTn+FaN/EYnmBqITd74aPc
0L+FemOybEQEMTqtMylPgok9KAtaIZcdCYaa3MCFCgw0dgL/gIIESt5zbx+/thgTaX78mVpIKpi6
heYMCsLefrDsEzjEaUyQ9zUK1Kodj1+9EmW0+5ksGuJtE5S2UzOig+CeJ420TL1yUXvz0srl8rKF
O6cx0WHejCoYZMwW/LFtR+oBikE6WwCDN+HYkgO6aXlM0QKsbv3dbD5QCoBIItVp1gS7qGhimUHD
Zp42oPxBxvphg7jljzT67KPLxT76RSBEFjD1foRtj+0tiR8D7d3Teq7kJyFH2+YrqgfaK1zkScPl
eEsvOGW4SGaRRUAGoY9U4XQlk4xU+JPadOQnUDJZGXIxM0IefbZbYxEis1TlKKCAaqRJNr7CryjT
UXvMqp0GucYR9gX7HFqICI6A38FE2wLopODBem3BUh6jSV8TBgg/adU6yFatqY3MEkKuvrksmFfE
1mqw1YUipHIKfPTYqJ4hYDbywWMYAv5Df7W7spd+8dgYejmyrZt11BAAxdoMjOSRTMDHPgcYR8lT
vCUo4x4+0T7zWmIMh29s5lc9MLn/+QMJAniVdJslC6mXrMi04fX+5p9VeSvjahluGyeiQ2KqT2kw
5RBx1LakdVqVokBhgduyoHkh19yE3smqbSw1CG/vQqcWW6CoEUJtnNEW9+Dm/EUik83dQRuzzhFu
MUZW92sgw+TzhXPc/ePCbEc+ETsiLIY/HLlpGjT8s8Q44iM9fQi+/+uigiSEV3f+Hout6XaSuoXc
ovdpS1wLfS1mtCC/LiRef+OExgQgVAIw+LMPPQiMilU4d1k5UFC/sD7Z4gw5UoqJmlL17QlkR+GE
RbKjmP1osHvtN4G2GFQu6HKDEUmhLmhSfvQCywut5HCBEeXTtIH4TrAZk8wCfZw2pNbjefYzJIXa
vIkAj/rygK6I8vJoNkeYmNHFlMkjWeDLSdDMP2z04QR0KrzxP987WH0kd9JMIA34pAmYARkuXQbw
6qrSMzLGFH7NtbMiZhdpJ8Qp+EkIx/vwGVNyEKAEnWQgukJB/PYND3nDLCaXZcdF686B0T8f06Jn
CPvF5lrNefmg6Mh1j0KbMhemmcfLYqmEl0KEFCHpj3TDQkkxeRta7u02Y8rzEoeI56A3FLlOL1u9
xHunGavTvhCbhxdjGZbLa7uq3e4F4H5kEOjEEbgG2n8YU96jDgR6gfxVoAx0EVVqyBA9luuFqDNW
OcpUvAij+pSIvt6zp2nqmJ3KodHeFyj8u3wu8x82GehDCHLgT2GSvSgY28v8nBemmb0/frW/pHwn
ah9NW+nvSXhmx0hkj++V84j8SeTm7FL0PYHZKMBZo2znXvQI9l1EY4xkuorjgMmxIvJW7NUVFHq9
6dNuxOVt/4WwNHb4sfHJORkzd63cDKyg2df3zSTtZQ1iDg+KbWYC6Cq25bLky7TLolJUunPPgGUx
0HGqyI0EAVCf6fr1D/USYCUsR4q+rOuX184DD8xpAsYiNwV8ad8imdAA9o0cvo0RLtga21SiW4FS
YS8sLZFK+apsUuS7nKMkJkj3fNZfOmhzW+9KiMUWegnpMHG1Bt/FUmPnPXeQSyRL4GlF2AH+bONw
M5KzxO4MmLhKS8NvwdNOwgyeR5/LM5OIj6PDN7AZn7S7YtijW0XUv1d833XOXnjxJqzQgRUr9UE6
cBcrSvmiQERhcUKP+d1kYqbrjsLiBSBDUI+pdQtVzSxzh4pVdGWjuu72RXO+6TMwtvJNoO8um2qk
jOGDAYYbFl/tBIe83lrfGpzOc2RxitqFiHn9ihiAeBr+Kb2haa/VCzOGT0JIv5PQg13R1xFVJGRt
I6itcAZ/GlnBydpA9Bt/4KSY/OlmdTgJgOfA5Onm3CAIq/HylhQLDRbV+kYQ4ux1BFZu04izlEQn
yCbs03NbMwZdUc8gfVCMFA2sFj6c8zjErOqJm6IYgq/Ze+nmYJjMVQ+dNg59g32xShtGUG/vEn7+
d1rALZKR96gPksyYYHkud0jRfIM1+5NP2nWfY3JflHfgqDj7IR35PrJYrtHRcyqtrfV45UVJcr53
v6XNxtJgyKM72aa8nC1FEpKCxQZwFvuGMV4XLoIODZ+VWkMv1CjsZ4rUvF8CeCmEiRd3EqOh0tIL
f09l1b3Bw+tzVdf2K6r3Zy8yaxOd3mW+eS5BbP4UcOMcVO6VeUli+AD9gVD2r4DUydXmiGy//cfP
mXlMTl3wlxDA09iArPoAg8CMQi9Nw5a1VJHRXf9kav5adD0V/MNEbw7r/V5QM+dM8sSS5uUzNwzL
cfzhx5hZEBmmAY8i/PvjKZnp+lwxX3OU/9XNDvDaMNJwEyOxVugwGyzR7TcjG+FxSmUzW+qYxS7W
WbIApF4HWY4VU2cMyn1cJz56okPZKjqLS+8IMKirl7mwNMuZsQ6j1NX7Ajl9EJKYU+SkJ4R0pvAl
NDHbheyghOwDiWjLL5VvcKMLQFcsb6xv1LkEh59mTIRbUc5UR+E2apluWyae6q4eZ1FX5lB0yeZM
2m6rdPSkZ3xrJchbG1ovoUtvs1zpvferLD3On9INdtU0KvsMGS2ivGmTetLTcIhjib16dmzBRC2j
WWQbAlL45Zd+OymW+6iHBlLVXOQYi6R2342F0u9pQw/49d9/R1WQWwkVidzWH8v7oNcBkG4IMMq7
TYI7xjK7C4GbdUBGOQG1B/GQ51a6sel6eh8Hlyc8KKbRhf1ZE4NWtKzXGLh+dbWhQEN0WGVSZhYr
hRbRkYng+xafdNukxthy0nr6OWM2j1GHaDmyRvyu2OZn0KxB78ZhIrZZ3SprvsfzqOlqXFXOg31k
kjB/RLF2QPtjDpxW2AIqtam3lc9zcnXboPiTjnVygOvCUm7y5famLUXTgGwQPIZhuL5GkBwqsR8L
qCsWK3dgq6+6tQfiV3qOwbhlx00AeZyfC7LAwdAT3hhMAHf2W5pZ/X3OwrHcjPU9GMsF4OusFM4K
6o3hPTH9eWqxi0xoZ1bPy086R5d/Hb5mBIwqheqmCqt3aMGoqSCPefaP3twmWWFmXq+JQILnGFp4
D03mXmlT7QVoPp+B9w9NNQ+gbnW3l3GH0Eb2C0JoYESUUCS2jiJ8wAm/LCNE97drwjxUfIgCHQDS
Pp0dL2WDjZwKAd9W7yZYCtxD5S2kggIa6XEEj+K8vBjtklKkhEbs3pPImdJtys3eIgt2i4Eb8Ihy
LcMgrlAFcpzshvsSlB1RXVDEYBhMQ+WZsyLlImI5nAziXT+8/1/nYexfDFBUEvCB9kBtLDx7nMby
tXCZPkwcPqmmsMhZ2T2s/jF8oUjFmbTBGHX3Dx3wqCXDGZ14xCqdsRk2SSnKO8GlY8H9U3byMHdi
p5EsoyezabUvgHWdwscmOPRW9jyzo0WmoVTlauTNYPeJLAs0fXdzSPnZGZp27eseqEdhpGTDtGv6
pknH0N9LKTNF0A1S7ENlNhDtWaRWxYd6UWOJ0+oNiNRuMgR4JRGKK54xotNXbhwKIcS9XTgeuInl
M3vKiVaKdKrBZAgNeYy7/3AQrcndpNgr+nkE6rwSKjyYM8XLEgY1dGl9Ypo/feJ+Igk3hwclr+NG
kJR60qDlHY4pdj3Vpy1K7JPZ6DHaoljDVOngpNporeN0/3jWbNVpaZivn60O/Jmozi20UTSQP3OE
RKvbDAvUymJSclIVfcbj9+mRdGlxtUjVqHcUNTqXYWWJbTp9wGlPh9zqAwOPvY7aaIfZq1MAZQlK
d1qYPTM9a7ehyDXpoonoELDMkrZVzccWdkI+tCs2CzSrofiXeWH1hgA+Lt65caf0IYcaG7QHJ0sh
a7ehFCzst1Etz8myl+ozi/6x8evBlHiADRTMYnue6WmuSD0cczC59YYzLy/Km6jQ9CbHo2hwl91V
lTHzvQbKJMhXn6LI8k1Is1SZjDbImIjkW3h0aV+5btOCOpJUzg9NG6ABXsePUz1r/J7T6+wQZmhu
Y5ycGv2csPNcatuOOCfQA8h9VeZcVybk1MLOBq2Al7lR0V/+udMNwJq+tFi4DFj53Byloa13U9dM
5a2F7Ex0iaxoT6WtYL2DOXx50wIbFTASu7sZMyuR0JR6cyXpUyi8lYg/UwO2IfJ+YQS4BxvYyUYn
sI05WVDAEKzkzqoA4QxS+5AovX3JdXZuTSxrfFTtByCff2U/pTkkIIaMBrgNIA9DAuFTvst7mGPE
DM6yOG65w8PtjSfSUOcwVnYsG4WoTxTxROTVnnq3ve2CXHMnfbFkpY0sauqoQThg6RPzEcunIvZn
TCVMAWOb1kT27fPu3JMzIWTdFrePSdFK3DJ9lCHOVoz4ZA2/9EGGw3OF9kL8lJdqdgUMxYhuSRWv
WWhWrdK2PriDeZUCiGenAfm7Akbp6y6VR0VWp+Lc3w9DhlC5gQSFrcS3sbXFfEmfhV6WgODWlYsZ
t0pP7zi7qF3EpSw6wd18wIOBNSOJAXckyuUrgia8xRIHQaSxWYTBIpV5zT6bKF69EZO6Xvg7rrSx
Wu7zuasgibLYsn7q6PXwFpLHLEX/PbYk4Zp/tL/4QADXkyGanKmenk/7fJ0d6OXcwNF2TCJ7Ll0t
Q5CF6wDeS5S7ayk5i27XvvZcWJVPDvJZ9LwtVmm5PbXp4KKlFt0gqXku4shAZ1xFxYdxpwr+P73S
o1kYxcgGejH6NP1PdkUB+n7mBXF9GCgOMs7+TPe8Imlri2ZHq+e0z2Oy3zLOWPwTALxPuyJMetP5
IIlGVmgwV7JG0RwKI7SETktbqZJAc5kGohA8sNCLHmxzINOIsd76sp7Gdidc034X0Do07XbDl+5H
BTM1SfGeQ3n6G5r0D9v8Yu9yTt/GpR74J8v2cdVsk73F0EaTE4zCo5+N4IZro4ly8ly837Ze2MB+
G940H8N8sknXlDXk6/AScfZIOquUMiBEO5w/2RxCkkJh6bGl7XtLNGTEPg59bw39gEkJjyyUW8ZG
O8HrXQ4a1aif7l7HIlbhR9GYGo/NQT9q8mF7Y78WYmjPGgL9qB67I3J3mRMzEEU/N4FLv1fAIhAh
f01NNGhLQObYpNKvKX83qMlkXBNJIQ5vdC4L7MnNnnfGmRjIiVS9vuUCnP75NFhBPYVTTd6gJGSH
IkmnaYX9ZbaA7/N9uEZcJWY2kWqsEGJKuZB4hvsa9S5HMP7eRyPhsq5qEa1qrHGdgxvliQ3fh6Tf
vFBJqOupaArHe6g6SXSOitU076GUhdTmFDIXmVRBvqy3Th2RDN3maFWYFuuJ1J8HQiTnq7Nux+aB
2rt6LG8NIsPIrXCVA+eY549Pi5HnolcLlKfqBJ/4QGVxWiZEQSZ2aefugDADA2vj1Qeo+mdQvuGM
VhJwfMPsKwVbjOwgny2EzoUD0/Dvu1YeUc8pay5ZYVA/80vNS6ptZlxPq59ohR5UpaA2EtoEcSDS
fChG69964u8CcHgF70OGzbMg5OgJO6MgWkeosZr6TE1rLtUr8B+TWY77aAwaHdFMd4ARdFzwuLZY
bg7ekmHjh87ryurjIm3nIfQJNgC5eV9gySojPoPRFS3Jqe+NBkoqT2lFYnMfXR4WyMtfH+BSyo5z
XMYqkXxq4QVJSxl70GyJeE6WWB2JOpO6I4cJwP+OdzazJhXnXVoj9nmIDoYKyQuzHclHrpCooOfU
59/5wHJebBDowS7HXhWkDUBrXuI67UGCfIYetrTS0qxAIwQwC2Zd6N3xFxHltqQ2AGUNLDWBKmNF
AXbl6edWMhkMBOK2cTQEeNzeLRsQW3vgkr7tRbxs4a+useSEcz7uv+YuJdtOEjEbSHmpn6Abe3rr
J+wSNDsG8zVYgVsfJJcJX1ufMJRlsV9TwggCaW8bPmvLd7VCynl+aaK23aKnc3mqgEHdgEoIgdUw
KpFLyimK3s2oHyAetejY+JnReeyGv/C0EFNzFegEWEHnPgfMLF/J2m9B6dyuAeP3H+8Qs8OB4Sir
t4I/mwJbXcNVCF2zY/Stqn2WaZLyxWDoHo3TqCPDpYyOsIRyn4fweYDh2fjm5+3ndkkwPKK61GP7
P+/yhZrHiwrl+rLq6nzeMDb1h1sEvSGgS5qgFPRss0ZIj3ZlSViHp5lECNq1t9v28cfjt4vPg7WG
QOD1JRIfFkW4RpNa89sf7JG86/0CS9ADwb10g5hvLhaUg7m19vZB5atVU2KTOuXmCcoP2rt/NFB6
XJwmhkXphMuoY9CUyMxoJ/U7mw+5nOBq2R2kslOT9rP8A5YP46o0PnSIjSUlxrZ5+8eY5NHeq7L4
s9hDUrxVX75Ua9sVEcpVNpR7MJOTv+JXO49fMYEHS3Az780BsEif+yg72MvzfA7Cny3xPq3jn0JB
cbu7xtbXaYYecDu9e61GgzKSHy1Twmb1/O+bqoVbohiomsvR+DisXxznrxwBc6AUjPnhhibBVn+K
Fq5Q1TiKS6nB2N8aA9aN+23xY5AX3MuX6BuJIRJg1SfVYiBnHGcOYcCg0RgEjsAHL2kT7IqvCFt0
qTlxuJuz4FcAaAZh0C7VNUOo+rEmLFiz7LJopLTPTRsFszZQ0Fwy3IAMwo+VmWsqJ4VJCLvEhBsJ
uNd8th+i4SSz7ne+xhbYEyA43BDsvr1wyYiLXUIAZmLsSyctimDFkEmE4bMS6yeHs51efYVVy1eg
qhCYwhI3nNz2w2vTEXHJBjkYRCDXJ98dFpAbBsSfNyx9eo1ItMLTBzkyT3T1Ew1+mm08HQNOHiOu
HP9EQEUplgbVRTqeHj4Lky/dCspOGtQNTpB8sMaxcj+Wje1XkZvzxYEoxTpH8T9U5rLrJLHGt8sP
x4zrv1iKkFGkoVDTm+5AGpxhyKrfljqFyYESnjnTaAWRhrG/soPkz6lCv7reJPmSNDpeWeu5zf5X
xiZZN87J2BVxtjork+phNejXFwqsItVS9Ek8WuKQpBF9WssZT5yITPrUrq96NvHEqwg++AcWKXV+
dlBsi/J8Ax4/fhBzTXBOsR3TYdKsy1swrRLYe6a/AAB05kvS+p2LD6Ofz9FObLzMqfIMT7C1LJe6
qRY8jyyH9DECKuncdsr5Bh/XlJ1UXcmTRcy50azi22X++yl4fA6QZz2gv2lASCJP5S9VqowMYNKc
kdl0FMuoh/IivNI0mlNrj2a9GIlFfG+om25whOtfZqrYN6i3kg4IAhwZDl4k2DPuRLKd4RY8/M4C
nSy8olImwtEVQrM1swJdavxqlQSB7iino1Yys+gKNTkWdQWGjQvS/Ewzz1yU1DC/6Mm3lxS62wRk
8SZFX302gqW7E7u0VxiFZMgStcrADT+TjeNaKvFVsCPMcQqn3OFtkbDJW3PEirlJ+TIasRRfSJRb
S5QIdfKhDZ4u37LmqK9FwXz1Losf0VbzQ6/SYsGpBqjYnUscMKF+Mjpsq9rgw44xnmzLK6H88SD1
FE60PPo65Mfm1fHNnsU5RQMP9Vr6WF8nB1WI2OvSdqKenEpL4SElfefhH9uxZN5uHNQ6LXQIXAoE
/XEERK5EQdRmYq4+fJcHxvItosH8dV75XPSxwCzN8w1pTXY6GnUqEsvADk6vZlz4LaR/5CjzqGS9
kjbnzNdTX+L+8CsiynmpPEFC3nDqe5FqGxHBPR5AGlPo90LLldvLOqvMBHu0ZCOD8mhUtQ9nK/1D
eev8du83X8rocCuE70sW3ie0N4t6n1/ryG4QO0z3g0TsQI4hl4+x4iA9q83yWeGQFhbhZZNX54sB
A9DhIy/ofTYCKnViiAa/y75RNCGnvGV7GMmmC7qi6YzCLLVLba7WkiToWgj5yfBQoLWpvfuDbeel
pfbHxVfuqBKkkUDiAQO7VA8tWyEyZBwtyYhUOgu+q1SQpxRkdeRISGyIm+ix+yqGOYoxqm/tBk5x
P8ETytsApgiSwGqXLUhGUjXHq3RThq96B65KLO4ZcHfzfrehwOUecBB0tPvxqXbxmrfkkQ4HbmSh
iorhen+UIW8fpFfEn9m5CVSFA0gUaDMNC55VDyMx1yFeCoYr826tviqJsfOv+6+W7fnWYQ6nqK+Z
azAlARB3Twz2ku4/gEhwmpwxH9Vqdjzbpa2TJSOeqlqOpqKfsKQ3/0AMCmM4TwI6G4GuO6UJw7UM
EseKm9IP2hK+TRIXjPtuWtNbFWITJopu46mdP1OQy0H/zSxf1cXbz6eSjTyjop5gMxjxzooCpB9s
xy3vjl+c3LNVrQ1OKwdE29qn3fwyZG7+gSvu0kRy3cWeczYoKNur9NcNqgIqkFsBq8D+y0DLGblq
sc5Vub5b1SMVYGEES5ZZlYyiSQpkfnCO0ftoMoYdVqbRFw+Yi8VrR9CQ2NFyG8UBChv3xPrr3hWw
ggnLQa6zPeR9XnwcksgLrlC0txo62gXej64GeAymVcQlQrhD7mKtwV/cPy7xAbHFs34hAUlasOAj
0O3rmA4/INLX2Vi6aDPbq9O6JfkVukuQ3jGl52fMGvczF5d4Y57v4+O9WVzMbDvBs2PGwAEzHLMp
YlNrNw2mX78/1s52yeKtAvctouL2oU4KiYU06Gm36hrtezM52+MQ4LeszM8XCBsYLuGySwJbTyJo
Co2ArC1o4VbYHIL3AyY6qywQY6kPRvDXclOBsf4eIJH9YFOwjppJGQgCbXNWjD/8kwCLhkvLFaNM
2w9XRWIB7oz4mEnWQZiIyb0TyVxWD46SRNfrXIt2s8YIMZXfAriFgWD1hmMAjNlvMP9o6TWcMaj5
JxW3+iBgTq4kxOZ/M3uCntbILGgTVNxrdhDWK9ViREMkD/RGpg765WhrrOSK59QzI4ZPb60nP2Qg
CO3/IuJriV/Mi8c/ctdl1ZbBkMljwGfPKhPjMLW5aKeFuKUx2ksH8ZT2r7NkOS/ZY7xwIvNWBL79
41SfNVPX7onjkhGG0N++yMdM9ewKEaTdtWEjjMVKM3z8kLTWXwh46qV6ssG9d5sfwCSxOOaFuogy
4/AEM1CrG2tIgk/KPd5CaPcRkGMUWanvrUJe4imbSjKbIXX89KEDzA1o308JnR3wW4Qw6ZE/0EUW
avf/vcFx/01BUcIMCXiATI6g6MAPvuuuIMdUEgbZacmtJpO0n6JaSzI6t07Ntim5kovy0BIVaG/8
dQQRUE2pQNqyk33UMi+W9Oi6oWto628Cla9udu/8uB45ypZlZCQhas1Dk1IY2QvdRtmIbfHk9oo7
9oQ7Qo90ghtUuSWMGQv6ztFCvgfNYP6bVbNQfl+w6qyeOCsybnmoXQAU3EBFdkymtgu44Y0WoNjr
TwIkmPtiYDgUhvuj3cRMlpvJ7NXy2EfIxjPkHFqtEEzAsJYwDVoRQ/8WcbTm4smcDM1u2jDd5py4
PE2sf6srcFPhLaA2RXAWSTkVxqvmQxWzsbQuqula95k/wTs2AayvwOr+Qwe4uvKcBwplmEUumyd7
AN+YtBjUv127ZmuBwOSbIKL6VO8fNXhPnjG3UpvLb/hxYyMETrmyn0FYgKTP0bOI5DF0ooUKRnbG
xta4sPbKkvMrZ/VU0rRjazwdhpNzX/u8iEehLH8nVvCSni7E6Rsa8nVGnXqGYJa5tSF78d9CkqGu
frkfu1fej7etwBbxijZLCrmmIANAYa72DVXYKUvvIJfD8r/OFV2ocB+cZtuJfGNTIjRd6CSxDMik
xLdYY09ZaBxH5WcMXbjFs3x4WyN3nd5tZAetUz7sazWvWcA=
`protect end_protected
